module Jvrki3(Yvrki3, Dwrki3, Lwrki3, Swrki3, Zwrki3, Jxrki3, Ayrki3, Lyrki3); 
`define L3lkc `AHB_DATA_WIDTH
parameter Xyrki3 = `L3lkc; 
input Yvrki3; 
input Dwrki3; 
input Lwrki3; 
input [(2 - 1):0] Swrki3; 
input Zwrki3; 
output Jxrki3; 
output [(2 - 1):0] Ayrki3; 
output [(Xyrki3 - 1):0] Lyrki3; 
reg Jxrki3; 
reg [(2 - 1):0] Ayrki3; 
reg Mzrki3; 
reg A0ski3; 
wire L0ski3; 
assign L0ski3 = (((Swrki3 == 2'b11) || (Swrki3 == 2'b10)) && ((Zwrki3 == 1'b1)  
&& (Lwrki3 == 1'b1))); 
assign Lyrki3 = {Xyrki3 {1'b0}}; 
always @(Mzrki3 or L0ski3) begin : Y0ski3 
case (Mzrki3) 
1'b0: begin 
if (L0ski3 == 1'b1) begin 
A0ski3 = 1'b1; 
end 
else begin 
A0ski3 = 1'b0; 
end 
end 
default: begin 
A0ski3 = 1'b0; 
end 
endcase 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : O1ski3 
if (Dwrki3 == 1'b0) begin 
Mzrki3 <= 1'b0; 
end 
else begin 
Mzrki3 <= A0ski3; 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : H2ski3 
if (Dwrki3 == 1'b0) begin 
Jxrki3 <= 1'b1; 
Ayrki3 <= 2'b0; 
end 
else 
begin 
case (Mzrki3) 
1'b0: begin 
if (L0ski3 == 1'b1) begin 
Jxrki3 <= 1'b0; 
Ayrki3 <= 2'b1; 
end 
else 
begin 
Jxrki3 <= 1'b1; 
Ayrki3 <= 2'b0; 
end 
end 
default: begin 
Jxrki3 <= 1'b1; 
Ayrki3 <= 2'b1; 
end 
endcase 
end 
end 
endmodule 
module R2ski3(Yvrki3, Dwrki3, D3ski3, J3ski3, U3ski3, H4ski3, S4ski3, F5ski3,  
Lwrki3, K5ski3, Q5ski3, U5ski3, B6ski3); 
input Yvrki3; 
input Dwrki3; 
input [(2 - 1):0] D3ski3; 
input [(32 - 1):0] J3ski3; 
input [(4 - 1):0] U3ski3; 
input F5ski3; 
input [3:0] H4ski3; 
input [((4 * 4) - 1):0] S4ski3; 
input Lwrki3; 
input Q5ski3; 
input K5ski3; 
output [(16 - 1):0] U5ski3; 
output [3:0] B6ski3; 
reg [(16 - 1):0] U5ski3; 
reg [3:0] B6ski3; 
reg [(32 - 1):0] G6ski3; 
reg [(16 - 1):0] T6ski3; 
reg E7ski3; 
reg [(2 - 1):0] Q7ski3; 
reg [3:0] C8ski3; 
reg [3:0] N8ski3; 
reg [(4 - 1):0] D9ski3; 
integer P9ski3; 
integer R9ski3; 
integer T9ski3; 
integer V9ski3; 
integer X9ski3; 
integer Z9ski3; 
integer Baski3; 
always @(J3ski3) begin : Daski3 
for (T9ski3 = 0; (T9ski3 <= (16 - 1)); T9ski3 = (T9ski3 + 1)) begin 
for (V9ski3 = 0; (V9ski3 < 2); V9ski3 = (V9ski3 + 1)) begin 
G6ski3[((T9ski3 * 2) + V9ski3)] = J3ski3[((16 * V9ski3) + T9ski3)]; 
end 
end 
end 
always @(G6ski3) begin : Uaski3 
U5ski3 = {16 {1'b0}}; 
for (X9ski3 = 0; (X9ski3 <= (16 - 1)); X9ski3 = (X9ski3 + 1)) begin 
Q7ski3 = (G6ski3 >> (2 * X9ski3)); 
U5ski3[X9ski3] = (|Q7ski3); 
end 
end 
always @(D3ski3 or T6ski3 or U5ski3 or U3ski3 or S4ski3 or F5ski3 or Lwrki3 or  
D9ski3 or H4ski3) begin : Gbski3 
B6ski3 = 16'b0; 
case (U3ski3) 
4'b1: 
Z9ski3 = 4; 
4'h2: 
Z9ski3 = 8; 
4'h3: 
Z9ski3 = 12; 
4'h4: 
Z9ski3 = 16; 
4'h5: 
Z9ski3 = 20; 
4'h6: 
Z9ski3 = 24; 
4'h7: 
Z9ski3 = 28; 
4'h8: 
Z9ski3 = 32; 
4'h9: 
Z9ski3 = 36; 
4'ha: 
Z9ski3 = 40; 
4'hb: 
Z9ski3 = 44; 
4'hc: 
Z9ski3 = 48; 
4'hd: 
Z9ski3 = 52; 
4'he: 
Z9ski3 = 56; 
4'hf: 
Z9ski3 = 60; 
default: 
Z9ski3 = 0; 
endcase 
N8ski3 = (S4ski3 >> Z9ski3); 
for (P9ski3 = 0; (P9ski3 < 4); P9ski3 = (P9ski3 + 1)) begin 
C8ski3 = (S4ski3 >> (4 * P9ski3)); 
B6ski3[P9ski3] = ((((((H4ski3[P9ski3] == 1'b1) || (D9ski3[P9ski3] == 1'b1)) || ( 
((D3ski3 == 2'b11) && (U3ski3 == P9ski3)) && (Lwrki3 == 1'b0))) || (( 
T6ski3[P9ski3] == 1'b1) && (U5ski3[P9ski3] == 1'b0))) || ((((F5ski3 == 1'b0) &&  
(D3ski3 == 2'b10)) && (C8ski3 > N8ski3)) && (Lwrki3 == 1'b0))) || ((((F5ski3 ==  
1'b1) && (D3ski3 == 2'b10)) && (U3ski3 != P9ski3)) && (Lwrki3 == 1'b0))); 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Qbski3 
if (Dwrki3 == 1'b0) begin 
T6ski3 <= {16 {1'b0}}; 
end 
else 
begin 
for (R9ski3 = 0; (R9ski3 < 16); R9ski3 = (R9ski3 + 1)) begin 
if (((D3ski3 == 2'b11) && (Lwrki3 == 1'b0)) && (U3ski3 == R9ski3)) begin 
T6ski3[R9ski3] <= 1'b1; 
end 
else 
begin 
if (U5ski3[R9ski3] == 1'b1) begin 
T6ski3[R9ski3] <= 1'b0; 
end 
end 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Gcski3 
if (Dwrki3 == 1'b0) begin 
E7ski3 <= {1'b0}; 
end 
else 
begin 
if (Lwrki3 == 1'b1) begin 
E7ski3 <= F5ski3; 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Xcski3 
if (Dwrki3 == 1'b0) begin 
D9ski3 <= {4 {1'b0}}; 
end 
else 
begin 
for (Baski3 = 0; (Baski3 < 4); Baski3 = (Baski3 + 1)) begin 
if (((((D3ski3 == 2'b11) && (E7ski3 == 1'b1)) && (Lwrki3 == 1'b0)) && (K5ski3 == 
1'b0)) && (U3ski3 != Baski3)) begin 
D9ski3[Baski3] <= 1'b1; 
end 
else 
begin 
if (Q5ski3 == 1'b1) begin 
D9ski3[Baski3] <= 1'b0; 
end 
end 
end 
end 
end 
endmodule 
module Odski3(Yvrki3, Dwrki3, Zdski3, Lwrki3, D3ski3, Keski3, Peski3, Veski3,  
Cfski3, Swrki3, Ifski3, Pfski3, Wfski3, Ggski3, J3ski3, U3ski3, Sgski3, Ygski3,  
Nhski3, Yhski3, Iiski3, Xiski3, Gjski3, Qjski3, Yjski3, Ikski3, Vkski3, Ilski3,  
Vlski3, Imski3, Vmski3, Inski3, Unski3, Goski3, Soski3, Epski3, Qpski3, Cqski3,  
Oqski3, Arski3, Mrski3, Yrski3); 
parameter Jsski3 = 32; 
parameter Xyrki3 = `L3lkc; 
`define M1lkc `BIG_ENDIAN
parameter Vsski3 = `M1lkc; 
input Yvrki3; 
input Dwrki3; 
input Zdski3; 
input Lwrki3; 
input [(2 - 1):0] D3ski3; 
input Keski3; 
input [(Jsski3 - 1):0] Peski3; 
input [(3 - 1):0] Veski3; 
input [(3 - 1):0] Cfski3; 
input [(2 - 1):0] Swrki3; 
input [(Xyrki3 - 1):0] Ifski3; 
input Pfski3; 
input [3:0] Wfski3; 
input [3:0] Ggski3; 
input [(32 - 1):0] J3ski3; 
input [(4 - 1):0] U3ski3; 
input Sgski3; 
input Ygski3; 
output [3:0] Nhski3; 
output Yhski3; 
output Iiski3; 
output [(2 - 1):0] Xiski3; 
output [(Xyrki3 - 1):0] Gjski3; 
output [(4 - 1):0] Qjski3; 
output Yjski3; 
output [(32 - 1):0] Ikski3; 
output [(32 - 1):0] Vkski3; 
output [(32 - 1):0] Ilski3; 
output [(32 - 1):0] Vlski3; 
output [(32 - 1):0] Imski3; 
output [(32 - 1):0] Vmski3; 
output [(32 - 1):0] Inski3; 
output [(32 - 1):0] Unski3; 
output [(32 - 1):0] Goski3; 
output [(32 - 1):0] Soski3; 
output [(32 - 1):0] Epski3; 
output [(32 - 1):0] Qpski3; 
output [(32 - 1):0] Cqski3; 
output [(32 - 1):0] Oqski3; 
output [(32 - 1):0] Arski3; 
output [3:1] Mrski3; 
output Yrski3; 
wire Gtski3; 
wire [((4 * 4) - 1):0] S4ski3; 
wire [(16 - 1):0] U5ski3; 
wire [9:0] Stski3; 
wire [(4 - 1):0] Buski3; 
wire [3:0] H4ski3; 
wire [3:0] B6ski3; 
wire [3:0] Juski3; 
wire [3:0] Tuski3; 
wire [3:0] Zuski3; 
wire [3:0] Ivski3; 
wire [3:0] Rvski3; 
wire Ewski3; 
wire Lwski3; 
wire Vwski3; 
wire Fxski3; 
wire Txski3; 
wire Zxski3; 
wire Kyski3; 
wire Syski3; 
wire Azski3; 
reg [255:0] Hzski3; 
wire Szski3; 
wire G0tki3; 
wire [3:0] S0tki3; 
wire [(480 - 1):0] F1tki3; 
wire R1tki3; 
wire [(32 - 1):0] W1tki3; 
wire Q5ski3; 
wire [(4 - 1):0] F2tki3; 
wire K5ski3; 
wire F5ski3; 
wire O2tki3; 
assign Mrski3[3:1] = ((0 == 1) ? Juski3[3:1] : {3 {1'b0}}); 
assign Yrski3 = ((0 == 1) ? Gtski3 : 1'b0); 
assign Kyski3 = ((1 == 0) ? 1'b0 : G0tki3); 
assign Yhski3 = ((1 == 0) ? 1'b0 : Szski3); 
assign Rvski3 = ((0 == 1'b1) ? Ivski3 : {3 {1'b0}}); 
assign Fxski3 = ((0 == 1'b1) ? Vwski3 : 1'b0); 
assign Qjski3 = F2tki3; 
C3tki3 #(Jsski3, Xyrki3, Vsski3) P3tki3( .Yvrki3 (Yvrki3),  .Dwrki3 (Dwrki3),  
.Keski3 (Keski3),  .Lwrki3 (Lwrki3),  .Qjski3 (F2tki3),  .Kyski3 (Kyski3),  
.Peski3 (Peski3),  .Swrki3 (Swrki3),  .Cfski3 (Cfski3),  .Ifski3 (Hzski3),  
.Pfski3 (Pfski3),  .Ygski3 (Ygski3),  .Iiski3 (Iiski3),  .Xiski3 (Xiski3),  
.Gjski3 (Gjski3),  .Zxski3 (Zxski3),  .Stski3 (Stski3),  .Txski3 (Txski3),  
.Buski3 (Buski3),  .S4ski3 (S4ski3),  .H4ski3 (H4ski3),  .R1tki3 (R1tki3),  
.F1tki3 (F1tki3),  .W1tki3 (W1tki3)); 
M4tki3 X4tki3( .Yvrki3 (Yvrki3),  .Dwrki3 (Dwrki3),  .Stski3 (Stski3),  .Txski3 
(Txski3),  .Zxski3 (Zxski3),  .Lwrki3 (Lwrki3),  .Syski3 (Syski3),  .O2tki3 
(O2tki3),  .F5ski3 (F5ski3),  .Yhski3 (Szski3),  .Kyski3 (G0tki3)); 
R2ski3 D5tki3( .Yvrki3 (Yvrki3),  .Dwrki3 (Dwrki3),  .D3ski3 (D3ski3),  .J3ski3 
(J3ski3),  .U3ski3 (U3ski3),  .H4ski3 (H4ski3),  .S4ski3 (S4ski3),  .F5ski3 
(F5ski3),  .K5ski3 (K5ski3),  .Lwrki3 (Lwrki3),  .Q5ski3 (Q5ski3),  .U5ski3 
(U5ski3),  .B6ski3 (B6ski3)); 
K5tki3 X5tki3( .Yvrki3 (Yvrki3),  .Dwrki3 (Dwrki3),  .Zdski3 (Zdski3),  .Wfski3 
(Wfski3),  .Buski3 (Buski3),  .Sgski3 (Sgski3),  .Veski3 (Veski3),  .Lwrki3 
(Lwrki3),  .D3ski3 (D3ski3),  .U5ski3 (U5ski3),  .Swrki3 (Swrki3),  .Zuski3 
(Zuski3),  .Lwski3 (Lwski3),  .B6ski3 (B6ski3),  .Kyski3 (Kyski3),  .Q5ski3 
(Q5ski3),  .O2tki3 (O2tki3),  .F5ski3 (F5ski3),  .K5ski3 (K5ski3),  .Ggski3 
(Ggski3),  .S0tki3 (S0tki3),  .Nhski3 (Nhski3),  .Yjski3 (Yjski3),  .Qjski3 
(F2tki3),  .Syski3 (Syski3)); 
F6tki3 #(4, 4, 1, 0, 0) T6tki3( .C7tki3 (Yvrki3),  .G7tki3 (Dwrki3),  .M7tki3 
(S0tki3),  .U7tki3 (S4ski3),  .D8tki3 ({(3 + 1) {1'b0}}),  .B6ski3 (B6ski3),  
.Ewski3 (Ewski3),  .Tuski3 (Tuski3)); 
C9tki3 Q9tki3( .R1tki3 (R1tki3),  .Zuski3 (Zuski3),  .Lwski3 (Lwski3),  .Tuski3 
(Tuski3),  .Ewski3 (Ewski3),  .Ivski3 (Rvski3),  .Vwski3 (Fxski3)); 
always @(Ifski3) begin : X3tki3 
Hzski3 = 256'b0; 
Hzski3[(Xyrki3 - 1):0] = Ifski3; 
end 
endmodule 
module M4tki3(Yvrki3, Dwrki3, Lwrki3, Stski3, Txski3, Zxski3, Syski3, F5ski3,  
O2tki3, Yhski3, Kyski3); 
parameter Z9tki3 = 2'b0; 
parameter Batki3 = 2'b1; 
parameter Datki3 = 2'b11; 
input Yvrki3; 
input Dwrki3; 
input Lwrki3; 
input [9:0] Stski3; 
input Txski3; 
input Zxski3; 
input Syski3; 
input F5ski3; 
input O2tki3; 
output Yhski3; 
output Kyski3; 
reg [9:0] Fatki3; 
wire [9:0] Patki3; 
reg Szski3; 
reg Vatki3; 
reg Ibtki3; 
wire Ybtki3; 
reg [1:0] Kctki3; 
wire [1:0] Mzrki3; 
reg [1:0] A0ski3; 
assign Mzrki3 = ((1 == 1'b1) ? Kctki3 : Z9tki3); 
assign Patki3 = ((1 == 1'b1) ? Fatki3 : 10'b0); 
assign Yhski3 = ((1 == 1'b1) ? Szski3 : 1'b0); 
assign Ybtki3 = ((1 == 1'b1) ? Ibtki3 : 1'b0); 
assign Kyski3 = (Vatki3 | Ybtki3); 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Cdtki3 
if (Dwrki3 == 1'b0) begin 
Kctki3 <= Z9tki3; 
end 
else begin 
Kctki3 <= A0ski3; 
end 
end 
always @(Mzrki3 or Txski3 or Syski3 or Patki3) begin : Y0ski3 
case (Mzrki3) 
Z9tki3: begin 
if ((Txski3 == 1'b1) && (Syski3 == 1'b1)) begin 
A0ski3 = Batki3; 
end 
else 
begin 
A0ski3 = Z9tki3; 
end 
end 
Batki3: begin 
if (Txski3 == 1'b1) begin 
if (Syski3 == 1'b1) begin 
A0ski3 = Batki3; 
end 
else 
begin 
if (Patki3 == 10'b1) begin 
A0ski3 = Datki3; 
end 
else 
begin 
A0ski3 = Batki3; 
end 
end 
end 
else 
begin 
A0ski3 = Z9tki3; 
end 
end 
Datki3: begin 
if (Txski3 == 1'b1) begin 
if (Syski3 == 1'b1) begin 
A0ski3 = Batki3; 
end 
else begin 
A0ski3 = Z9tki3; 
end 
end 
else 
begin 
A0ski3 = Z9tki3; 
end 
end 
default: 
A0ski3 = Z9tki3; 
endcase 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Udtki3 
if (Dwrki3 == 1'b0) begin 
Fatki3 <= 10'b0; 
end 
else 
begin 
if (Mzrki3 == Datki3) begin 
Fatki3 <= Stski3; 
end 
else 
begin 
if (Syski3 == 1'b1) begin 
Fatki3 <= Stski3; 
end 
else 
begin 
if (Fatki3 == 10'b0) begin 
Fatki3 <= Fatki3; 
end 
else 
begin 
Fatki3 <= (Fatki3 - 10'b1); 
end 
end 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Fetki3 
if (Dwrki3 == 1'b0) begin 
Szski3 <= 1'b0; 
end 
else 
begin 
if (Txski3 == 1'b0) begin 
Szski3 <= 1'b0; 
end 
else 
begin 
if ((((Kyski3 == 1'b1) && (Lwrki3 == 1'b1)) && (F5ski3 == 1'b0)) && (O2tki3 ==  
1'b0)) begin 
Szski3 <= 1'b1; 
end 
else 
begin 
if (Zxski3 == 1'b1) begin 
Szski3 <= 1'b0; 
end 
end 
end 
end 
end 
always @(Mzrki3 or Txski3) begin : Uetki3 
if (Mzrki3 == Datki3) begin 
Vatki3 = Txski3; 
end 
else 
begin 
Vatki3 = 1'b0; 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Mftki3 
if (Dwrki3 == 1'b0) begin 
Ibtki3 <= 1'b0; 
end 
else 
begin 
if (Txski3 == 1'b1) begin 
if (Lwrki3 == 1'b0) begin 
if (Vatki3 == 1'b1) begin 
Ibtki3 <= 1'b1; 
end 
end 
else 
begin 
Ibtki3 <= 1'b0; 
end 
end 
else 
begin 
Ibtki3 <= 1'b0; 
end 
end 
end 
endmodule 
module Dgtki3(Yvrki3, Dwrki3, Ogtki3, Ygtki3, Qjski3, Jhtki3, Thtki3, Ditki3,  
Oitki3, Zitki3, Lyrki3, Jxrki3, Ayrki3, Kjtki3, Vjtki3, Fktki3, Keski3, U3ski3,  
Peski3, Veski3, Qktki3, Cfski3, Swrki3, Ifski3, Pfski3, Wktki3, Lwrki3, D3ski3); 
parameter Jsski3 = 32; 
parameter Xyrki3 = `L3lkc; 
parameter Dltki3 = ((3 + 1) * Jsski3); 
parameter Rltki3 = (4 * Xyrki3); 
parameter Fmtki3 = (3 * Xyrki3); 
input Yvrki3; 
input Dwrki3; 
input [(Dltki3 - 1):0] Ogtki3; 
input [(12 - 1):0] Ygtki3; 
input [(4 - 1):0] Qjski3; 
input [(16 - 1):0] Jhtki3; 
input [(12 - 1):0] Thtki3; 
input [(8 - 1):0] Ditki3; 
input [(Rltki3 - 1):0] Oitki3; 
input [(4 - 1):0] Zitki3; 
input [(Xyrki3 - 1):0] Lyrki3; 
input [(Fmtki3 - 1):0] Fktki3; 
input Jxrki3; 
input [(2 - 1):0] Ayrki3; 
input [(3 - 1):0] Kjtki3; 
input [(6 - 1):0] Vjtki3; 
input [2:0] Keski3; 
output [(Jsski3 - 1):0] Peski3; 
output [(3 - 1):0] Veski3; 
output [(4 - 1):0] Qktki3; 
output [(3 - 1):0] Cfski3; 
output [(2 - 1):0] Swrki3; 
output [(Xyrki3 - 1):0] Ifski3; 
output Pfski3; 
output [(4 - 1):0] U3ski3; 
output [(Xyrki3 - 1):0] Wktki3; 
output Lwrki3; 
output [(2 - 1):0] D3ski3; 
reg [(Xyrki3 - 1):0] Wktki3; 
reg Lwrki3; 
reg [(2 - 1):0] D3ski3; 
reg [(4 - 1):0] Vmtki3; 
wire [(4 - 1):0] F2tki3; 
reg [2:0] Jntki3; 
integer R9ski3; 
assign U3ski3 = ((0 == 1'b1) ? 4'b1 : Vmtki3); 
assign F2tki3 = ((0 == 1'b1) ? 4'b1 : Qjski3); 
Tntki3 #(Dltki3, 4, Jsski3) Gotki3( .Kotki3 (Ogtki3),  .Motki3 (F2tki3),  
.Qotki3 (Peski3)); 
Tntki3 #(8, 4, 2) Uotki3( .Kotki3 (Ditki3),  .Motki3 (F2tki3),  .Qotki3 (Swrki3) 
); 
Tntki3 #(12, 4, 3) Yotki3( .Kotki3 (Ygtki3),  .Motki3 (F2tki3),  .Qotki3 
(Veski3)); 
Tntki3 #(12, 4, 3) Cptki3( .Kotki3 (Thtki3),  .Motki3 (F2tki3),  .Qotki3 
(Cfski3)); 
Tntki3 #(16, 4, 4) Gptki3( .Kotki3 (Jhtki3),  .Motki3 (F2tki3),  .Qotki3 
(Qktki3)); 
Tntki3 #(4, 4, 1) Kptki3( .Kotki3 (Zitki3),  .Motki3 (F2tki3),  .Qotki3 (Pfski3) 
); 
Tntki3 #(Rltki3, 4, Xyrki3) Pptki3( .Kotki3 (Oitki3),  .Motki3 (U3ski3),  
.Qotki3 (Ifski3)); 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Uptki3 
if (Dwrki3 == 1'b0) begin 
Vmtki3 <= {4 {1'b0}}; 
end 
else 
begin 
if (Lwrki3 == 1'b1) begin 
Vmtki3 <= Qjski3; 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Mqtki3 
if (Dwrki3 == 1'b0) begin 
Jntki3 <= {(2 + 1) {1'b0}}; 
end 
else 
begin 
if (Lwrki3 == 1'b1) begin 
if (Swrki3 == 2'b0) begin 
Jntki3 <= {(2 + 1) {1'b0}}; 
end 
else 
begin 
Jntki3 <= Keski3; 
end 
end 
end 
end 
always @(Jntki3 or Fktki3 or Kjtki3 or Vjtki3 or Ayrki3 or Lyrki3 or Jxrki3)  
begin : Brtki3 
Lwrki3 = Jxrki3; 
D3ski3 = Ayrki3; 
Wktki3 = Lyrki3; 
for (R9ski3 = 0; (R9ski3 <= 2); R9ski3 = (R9ski3 + 1)) begin 
if (Jntki3[R9ski3] == 1'b1) begin 
Lwrki3 = Kjtki3[R9ski3]; 
D3ski3 = (Vjtki3 >> (R9ski3 * 2)); 
Wktki3 = (Fktki3 >> (R9ski3 * Xyrki3)); 
end 
end 
end 
endmodule 
module C3tki3(Yvrki3, Dwrki3, Keski3, Lwrki3, Qjski3, Kyski3, Peski3, Swrki3,  
Cfski3, Ifski3, Pfski3, Ygski3, Iiski3, Xiski3, Gjski3, Zxski3, Stski3, Txski3,  
Buski3, S4ski3, H4ski3, R1tki3, F1tki3, W1tki3); 
parameter Jsski3 = 32; 
parameter Xyrki3 = `L3lkc; 
parameter Vsski3 = `M1lkc; 
parameter O9uki3 = 2'b0; 
parameter W9uki3 = 2'b1; 
parameter Eauki3 = 2'b10; 
parameter Nauki3 = 2'b11; 
input Yvrki3; 
input Dwrki3; 
input Keski3; 
input Lwrki3; 
input [(4 - 1):0] Qjski3; 
input Kyski3; 
input [(Jsski3 - 1):0] Peski3; 
input [(2 - 1):0] Swrki3; 
input [(3 - 1):0] Cfski3; 
input [255:0] Ifski3; 
input Pfski3; 
input Ygski3; 
output Iiski3; 
output [(2 - 1):0] Xiski3; 
output [(Xyrki3 - 1):0] Gjski3; 
output [9:0] Stski3; 
output Txski3; 
output [(4 - 1):0] Buski3; 
output Zxski3; 
output [((4 * 4) - 1):0] S4ski3; 
output [3:0] H4ski3; 
output R1tki3; 
output [(480 - 1):0] F1tki3; 
output [(32 - 1):0] W1tki3; 
reg Zxski3; 
wire L0ski3; 
wire Xrtki3; 
wire Hstki3; 
wire Rstki3; 
wire Zstki3; 
wire Httki3; 
wire Pttki3; 
wire Xttki3; 
wire Futki3; 
wire Nutki3; 
wire Vutki3; 
wire Dvtki3; 
wire Lvtki3; 
wire Uvtki3; 
wire Dwtki3; 
wire Mwtki3; 
wire Vwtki3; 
wire Extki3; 
wire Nxtki3; 
wire Aytki3; 
wire Kytki3; 
wire Wytki3; 
wire [255:0] Aztki3; 
wire [15:0] Oztki3; 
wire [63:0] D0uki3; 
wire [3:0] U0uki3; 
wire [3:0] E1uki3; 
wire [3:0] O1uki3; 
wire [3:0] Y1uki3; 
wire [3:0] I2uki3; 
wire [3:0] S2uki3; 
wire [3:0] C3uki3; 
wire [3:0] M3uki3; 
wire [3:0] W3uki3; 
wire [3:0] G4uki3; 
wire [3:0] R4uki3; 
wire [3:0] C5uki3; 
wire [3:0] N5uki3; 
wire [3:0] Y5uki3; 
wire [3:0] J6uki3; 
wire [9:0] U6uki3; 
wire [9:0] E7uki3; 
wire [(4 - 1):0] T7uki3; 
wire G8uki3; 
wire Q8uki3; 
wire C9uki3; 
reg [3:0] Wauki3; 
reg [3:0] Bbuki3; 
reg [3:0] Gbuki3; 
reg [3:0] Lbuki3; 
reg [3:0] Qbuki3; 
reg [3:0] Vbuki3; 
reg [3:0] Acuki3; 
reg [3:0] Fcuki3; 
reg [3:0] Kcuki3; 
reg [3:0] Pcuki3; 
reg [3:0] Vcuki3; 
reg [3:0] Bduki3; 
reg [3:0] Hduki3; 
reg [3:0] Nduki3; 
reg [3:0] Tduki3; 
wire [3:0] Zduki3; 
wire [3:0] Deuki3; 
wire [3:0] Heuki3; 
wire [3:0] Leuki3; 
wire [3:0] Peuki3; 
wire [3:0] Teuki3; 
wire [3:0] Xeuki3; 
wire [3:0] Bfuki3; 
wire [3:0] Ffuki3; 
wire [3:0] Jfuki3; 
wire [3:0] Ofuki3; 
wire [3:0] Tfuki3; 
wire [3:0] Yfuki3; 
wire [3:0] Dguki3; 
wire [3:0] Iguki3; 
reg [9:0] Nguki3; 
reg Xguki3; 
reg [3:0] Ehuki3; 
reg Nhuki3; 
reg Eiuki3; 
reg [(2 - 1):0] Uiuki3; 
reg Fjuki3; 
reg Qjuki3; 
reg [(4 - 1):0] Dkuki3; 
reg [(Jsski3 - 1):0] Pkuki3; 
reg [(2 - 1):0] Zkuki3; 
reg [(3 - 1):0] Kluki3; 
wire [(Jsski3 - 1):0] Uluki3; 
wire [(2 - 1):0] Cmuki3; 
wire [(3 - 1):0] Lmuki3; 
wire Tmuki3; 
wire Cnuki3; 
wire [(4 - 1):0] Nnuki3; 
reg [1:0] Xnuki3; 
wire [1:0] Fouki3; 
reg [1:0] Louki3; 
reg [31:0] Vouki3; 
reg [31:0] Gpuki3; 
reg [31:0] Opuki3; 
reg Aquki3; 
wire Iquki3; 
reg Mquki3; 
wire [(32 - 1):0] Yquki3; 
wire [(32 - 1):0] Nruki3; 
wire [(32 - 1):0] Csuki3; 
wire [(32 - 1):0] Rsuki3; 
wire [(32 - 1):0] Gtuki3; 
wire [(32 - 1):0] Vtuki3; 
wire [(32 - 1):0] Kuuki3; 
wire [(32 - 1):0] Zuuki3; 
wire [(32 - 1):0] Ovuki3; 
wire [(32 - 1):0] Dwuki3; 
wire [(32 - 1):0] Twuki3; 
wire [(32 - 1):0] Jxuki3; 
wire [(32 - 1):0] Zxuki3; 
wire [(32 - 1):0] Pyuki3; 
wire [(32 - 1):0] Fzuki3; 
reg Vzuki3; 
wire B0vki3; 
wire M0vki3; 
reg [31:0] V0vki3; 
reg [31:0] L1vki3; 
reg [31:0] B2vki3; 
reg [31:0] R2vki3; 
reg [31:0] H3vki3; 
reg [31:0] X3vki3; 
reg [31:0] N4vki3; 
reg [31:0] D5vki3; 
reg [31:0] T5vki3; 
reg [31:0] J6vki3; 
reg [31:0] A7vki3; 
reg [31:0] R7vki3; 
reg [31:0] I8vki3; 
reg [31:0] Z8vki3; 
reg [31:0] Q9vki3; 
wire [(32 - 1):0] Havki3; 
wire [(32 - 1):0] Vavki3; 
reg [(32 - 1):0] Fbvki3; 
reg [31:0] Obvki3; 
wire Acvki3; 
reg [(32 - 1):0] Mcvki3; 
reg [(32 - 1):0] Ycvki3; 
reg [(32 - 1):0] Kdvki3; 
reg [(32 - 1):0] Wdvki3; 
reg [(32 - 1):0] Ievki3; 
reg [(32 - 1):0] Uevki3; 
reg [(32 - 1):0] Gfvki3; 
reg [(32 - 1):0] Sfvki3; 
reg [(32 - 1):0] Egvki3; 
reg [(32 - 1):0] Qgvki3; 
reg [(32 - 1):0] Dhvki3; 
reg [(32 - 1):0] Qhvki3; 
reg [(32 - 1):0] Divki3; 
reg [(32 - 1):0] Qivki3; 
reg [(32 - 1):0] Djvki3; 
wire [(32 - 1):0] Qjvki3; 
wire [(32 - 1):0] Dkvki3; 
wire [(32 - 1):0] Qkvki3; 
wire [(32 - 1):0] Dlvki3; 
wire [(32 - 1):0] Qlvki3; 
wire [(32 - 1):0] Dmvki3; 
wire [(32 - 1):0] Qmvki3; 
wire [(32 - 1):0] Dnvki3; 
wire [(32 - 1):0] Qnvki3; 
wire [(32 - 1):0] Dovki3; 
wire [(32 - 1):0] Rovki3; 
wire [(32 - 1):0] Fpvki3; 
wire [(32 - 1):0] Tpvki3; 
wire [(32 - 1):0] Hqvki3; 
wire [(32 - 1):0] Vqvki3; 
wire [(32 - 1):0] Jrvki3; 
wire [(32 - 1):0] Asvki3; 
wire [(32 - 1):0] Rsvki3; 
wire [(32 - 1):0] Itvki3; 
wire [(32 - 1):0] Ztvki3; 
wire [(32 - 1):0] Quvki3; 
wire [(32 - 1):0] Hvvki3; 
wire [(32 - 1):0] Yvvki3; 
wire [(32 - 1):0] Pwvki3; 
wire [(32 - 1):0] Gxvki3; 
wire [(32 - 1):0] Yxvki3; 
wire [(32 - 1):0] Qyvki3; 
wire [(32 - 1):0] Izvki3; 
wire [(32 - 1):0] A0wki3; 
wire [(32 - 1):0] S0wki3; 
wire K1wki3; 
wire V1wki3; 
wire G2wki3; 
wire R2wki3; 
wire C3wki3; 
wire N3wki3; 
wire Y3wki3; 
wire J4wki3; 
wire U4wki3; 
wire F5wki3; 
wire R5wki3; 
wire D6wki3; 
wire P6wki3; 
wire B7wki3; 
wire N7wki3; 
wire Z7wki3; 
wire [31:0] R8wki3; 
assign L0ski3 = ((Swrki3 != 2'b0) && (Swrki3 != 2'b1)); 
assign Xrtki3 = ((Keski3 == 1'b1) && (Lwrki3 == 1'b1)); 
assign Hstki3 = ((Xrtki3 == 1'b1) && (L0ski3 == 1'b1)); 
assign Cnuki3 = ((1 == 1) ? Qjuki3 : 1'b0); 
assign Tmuki3 = ((1 == 1) ? Fjuki3 : 1'b0); 
assign Uluki3 = ((1 == 1) ? Pkuki3 : {Jsski3 {1'b0}}); 
assign Cmuki3 = ((1 == 1) ? Zkuki3 : {2 {1'b0}}); 
assign Lmuki3 = ((1 == 1) ? Kluki3 : {4 {1'b0}}); 
assign Nnuki3 = ((1 == 1) ? Dkuki3 : {4 {1'b0}}); 
assign G8uki3 = ((Cmuki3 != 2'b0) && (Cmuki3 != 2'b1)); 
assign Q8uki3 = ((G8uki3 == 1'b1) && (Cnuki3 == 1'b1)); 
assign Xiski3 = ((1 == 1'b1) ? Uiuki3 : {2 {1'b0}}); 
assign Iiski3 = ((1 == 1'b1) ? Nhuki3 : 1'b1); 
assign Fouki3 = ((1 == 1'b1) ? Xnuki3 : O9uki3); 
assign Wytki3 = (((Tmuki3 == 1'b1) && (Q8uki3 == 1'b1)) && (Lwrki3 == 1'b1)); 
assign Rstki3 = ((Uluki3[9:0] == 10'b0) && (Wytki3 == 1'b1)); 
assign Zstki3 = ((Uluki3[9:0] == 10'h004) && (Wytki3 == 1'b1)); 
assign Httki3 = ((Uluki3[9:0] == 10'h008) && (Wytki3 == 1'b1)); 
assign Pttki3 = ((Uluki3[9:0] == 10'h00c) && (Wytki3 == 1'b1)); 
assign Xttki3 = ((Uluki3[9:0] == 10'h010) && (Wytki3 == 1'b1)); 
assign Futki3 = ((Uluki3[9:0] == 10'h014) && (Wytki3 == 1'b1)); 
assign Nutki3 = ((Uluki3[9:0] == 10'h018) && (Wytki3 == 1'b1)); 
assign Vutki3 = ((Uluki3[9:0] == 10'h01c) && (Wytki3 == 1'b1)); 
assign Dvtki3 = ((Uluki3[9:0] == 10'h020) && (Wytki3 == 1'b1)); 
assign Lvtki3 = ((Uluki3[9:0] == 10'h024) && (Wytki3 == 1'b1)); 
assign Uvtki3 = ((Uluki3[9:0] == 10'h028) && (Wytki3 == 1'b1)); 
assign Dwtki3 = ((Uluki3[9:0] == 10'h02c) && (Wytki3 == 1'b1)); 
assign Mwtki3 = ((Uluki3[9:0] == 10'h030) && (Wytki3 == 1'b1)); 
assign Vwtki3 = ((Uluki3[9:0] == 10'h034) && (Wytki3 == 1'b1)); 
assign Extki3 = ((Uluki3[9:0] == 10'h038) && (Wytki3 == 1'b1)); 
assign Nxtki3 = ((Uluki3[9:0] == 10'h03c) && (Wytki3 == 1'b1)); 
assign Aytki3 = ((Uluki3[9:0] == 10'h040) && (Wytki3 == 1'b1)); 
assign Kytki3 = ((Uluki3[9:0] == 10'h048) && (Wytki3 == 1'b1)); 
assign M0vki3 = ((Uluki3[9:0] == 10'h04c) && (Wytki3 == 1'b1)); 
assign Acvki3 = ((Uluki3[9:0] == 10'h050) && (Wytki3 == 1'b1)); 
assign K1wki3 = ((Uluki3[9:0] == 10'h054) && (Wytki3 == 1'b1)); 
assign V1wki3 = ((Uluki3[9:0] == 10'h058) && (Wytki3 == 1'b1)); 
assign G2wki3 = ((Uluki3[9:0] == 10'h05c) && (Wytki3 == 1'b1)); 
assign R2wki3 = ((Uluki3[9:0] == 10'h060) && (Wytki3 == 1'b1)); 
assign C3wki3 = ((Uluki3[9:0] == 10'h064) && (Wytki3 == 1'b1)); 
assign N3wki3 = ((Uluki3[9:0] == 10'h068) && (Wytki3 == 1'b1)); 
assign Y3wki3 = ((Uluki3[9:0] == 10'h06c) && (Wytki3 == 1'b1)); 
assign J4wki3 = ((Uluki3[9:0] == 10'h070) && (Wytki3 == 1'b1)); 
assign U4wki3 = ((Uluki3[9:0] == 10'h074) && (Wytki3 == 1'b1)); 
assign F5wki3 = ((Uluki3[9:0] == 10'h078) && (Wytki3 == 1'b1)); 
assign R5wki3 = ((Uluki3[9:0] == 10'h07c) && (Wytki3 == 1'b1)); 
assign D6wki3 = ((Uluki3[9:0] == 10'h080) && (Wytki3 == 1'b1)); 
assign P6wki3 = ((Uluki3[9:0] == 10'h084) && (Wytki3 == 1'b1)); 
assign B7wki3 = ((Uluki3[9:0] == 10'h088) && (Wytki3 == 1'b1)); 
assign N7wki3 = ((Uluki3[9:0] == 10'h08c) && (Wytki3 == 1'b1)); 
assign Z7wki3 = ((0 == 1'b1) ? (Ygski3 == 1'b0) : (Vsski3 == 1'b0)); 
assign U0uki3 = Vouki3[3:0]; 
assign Zduki3 = (((1 == 0) || (0 == 1)) ? 4'b1 : Wauki3); 
assign E1uki3 = Vouki3[3:0]; 
assign Deuki3 = ((3 < 2) ? 4'b0 : (((1 == 0) || (0 == 1)) ? 4'h2 : Bbuki3)); 
assign O1uki3 = Vouki3[3:0]; 
assign Heuki3 = ((3 < 3) ? 4'b0 : (((1 == 0) || (0 == 1)) ? 4'h3 : Gbuki3)); 
assign Y1uki3 = Vouki3[3:0]; 
assign Leuki3 = ((3 < 4) ? 4'b0 : (((1 == 0) || (0 == 1)) ? 4'h4 : Lbuki3)); 
assign I2uki3 = Vouki3[3:0]; 
assign Peuki3 = ((3 < 5) ? 4'b0 : (((1 == 0) || (0 == 1)) ? 4'h5 : Qbuki3)); 
assign S2uki3 = Vouki3[3:0]; 
assign Teuki3 = ((3 < 6) ? 4'b0 : (((1 == 0) || (0 == 1)) ? 4'h6 : Vbuki3)); 
assign C3uki3 = Vouki3[3:0]; 
assign Xeuki3 = ((3 < 7) ? 4'b0 : (((1 == 0) || (0 == 1)) ? 4'h7 : Acuki3)); 
assign M3uki3 = Vouki3[3:0]; 
assign Bfuki3 = ((3 < 8) ? 4'b0 : (((1 == 0) || (0 == 1)) ? 4'h8 : Fcuki3)); 
assign W3uki3 = Vouki3[3:0]; 
assign Ffuki3 = ((3 < 9) ? 4'b0 : (((1 == 0) || (0 == 1)) ? 4'h9 : Kcuki3)); 
assign G4uki3 = Vouki3[3:0]; 
assign Jfuki3 = ((3 < 10) ? 4'b0 : (((1 == 0) || (0 == 1)) ? 4'ha : Pcuki3)); 
assign R4uki3 = Vouki3[3:0]; 
assign Ofuki3 = ((3 < 11) ? 4'b0 : (((1 == 0) || (0 == 1)) ? 4'hb : Vcuki3)); 
assign C5uki3 = Vouki3[3:0]; 
assign Tfuki3 = ((3 < 12) ? 4'b0 : (((1 == 0) || (0 == 1)) ? 4'hc : Bduki3)); 
assign N5uki3 = Vouki3[3:0]; 
assign Yfuki3 = ((3 < 13) ? 4'b0 : (((1 == 0) || (0 == 1)) ? 4'hd : Hduki3)); 
assign Y5uki3 = Vouki3[3:0]; 
assign Dguki3 = ((3 < 14) ? 4'b0 : (((1 == 0) || (0 == 1)) ? 4'he : Nduki3)); 
assign J6uki3 = Vouki3[3:0]; 
assign Iguki3 = ((3 < 15) ? 4'b0 : (((1 == 0) || (0 == 1)) ? 4'hf : Tduki3)); 
assign E7uki3 = Vouki3[9:0]; 
assign C9uki3 = Vouki3[0]; 
assign Stski3 = (((1 == 1'b0) || (1 == 1'b0)) ? 10'b0 : Nguki3); 
assign Txski3 = (((1 == 1'b0) || (1 == 1'b0)) ? 1'b0 : Xguki3); 
assign T7uki3 = Vouki3[3:0]; 
assign Buski3 = (((0 == 1) || (1 == 1'b0)) ? 0 : Ehuki3); 
assign Iquki3 = (((1 == 1'b1) && (1 == 1'b1)) ? Aquki3 : 1'b0); 
assign B0vki3 = Vouki3[0]; 
assign R1tki3 = (((0 == 1'b1) && (1 == 1'b1)) ? Vzuki3 : 1'b0); 
assign Havki3 = Vouki3[(32 - 1):0]; 
assign Vavki3 = (((1 == 1) || (1 == 1'b0)) ? 32'h0000ffff : Fbvki3); 
assign W1tki3 = Vavki3; 
assign Jrvki3 = Vouki3[(32 - 1):0]; 
assign Qjvki3 = (((1 == 1) || (1 == 1'b0)) ? 32'h0000000f : Mcvki3); 
assign Asvki3 = Vouki3[(32 - 1):0]; 
assign Dkvki3 = (((1 == 1) || (1 == 1'b0)) ? 32'h0000000f : Ycvki3); 
assign Rsvki3 = Vouki3[(32 - 1):0]; 
assign Qkvki3 = (((1 == 1) || (1 == 1'b0)) ? 32'h0000000f : Kdvki3); 
assign Itvki3 = Vouki3[(32 - 1):0]; 
assign Dlvki3 = (((1 == 1) || (1 == 1'b0)) ? 32'h0000000f : Wdvki3); 
assign Ztvki3 = Vouki3[(32 - 1):0]; 
assign Qlvki3 = (((1 == 1) || (1 == 1'b0)) ? 32'h0000000f : Ievki3); 
assign Quvki3 = Vouki3[(32 - 1):0]; 
assign Dmvki3 = (((1 == 1) || (1 == 1'b0)) ? 32'h0000000f : Uevki3); 
assign Hvvki3 = Vouki3[(32 - 1):0]; 
assign Qmvki3 = (((1 == 1) || (1 == 1'b0)) ? 32'h0000000f : Gfvki3); 
assign Yvvki3 = Vouki3[(32 - 1):0]; 
assign Dnvki3 = (((1 == 1) || (1 == 1'b0)) ? 32'h0000000f : Sfvki3); 
assign Pwvki3 = Vouki3[(32 - 1):0]; 
assign Qnvki3 = (((1 == 1) || (1 == 1'b0)) ? 32'h0000000f : Egvki3); 
assign Gxvki3 = Vouki3[(32 - 1):0]; 
assign Dovki3 = (((1 == 1) || (1 == 1'b0)) ? 32'h0000000f : Qgvki3); 
assign Yxvki3 = Vouki3[(32 - 1):0]; 
assign Rovki3 = (((1 == 1) || (1 == 1'b0)) ? 32'h0000000f : Dhvki3); 
assign Qyvki3 = Vouki3[(32 - 1):0]; 
assign Fpvki3 = (((1 == 1) || (1 == 1'b0)) ? 32'h0000000f : Qhvki3); 
assign Izvki3 = Vouki3[(32 - 1):0]; 
assign Tpvki3 = (((1 == 1) || (1 == 1'b0)) ? 32'h0000000f : Divki3); 
assign A0wki3 = Vouki3[(32 - 1):0]; 
assign Hqvki3 = (((1 == 1) || (1 == 1'b0)) ? 32'h0000000f : Qivki3); 
assign S0wki3 = Vouki3[(32 - 1):0]; 
assign Vqvki3 = (((1 == 1) || (1 == 1'b0)) ? 32'h0000000f : Djvki3); 
assign U6uki3 = (Iiski3 ? Peski3[9:0] : Uluki3[9:0]); 
assign R8wki3 = 32'h3230312a; 
assign Aztki3[31:0] = ((Z7wki3 == 1'b1) ? Gpuki3[31:0] : {Gpuki3[7:0],  
Gpuki3[15:8], Gpuki3[23:16], Gpuki3[31:24]}); 
assign Aztki3[63:32] = Aztki3[31:0]; 
assign Aztki3[95:64] = Aztki3[31:0]; 
assign Aztki3[127:96] = Aztki3[31:0]; 
assign Aztki3[159:128] = Aztki3[31:0]; 
assign Aztki3[191:160] = Aztki3[31:0]; 
assign Aztki3[223:192] = Aztki3[31:0]; 
assign Aztki3[255:224] = Aztki3[31:0]; 
assign Gjski3 = Aztki3[(Xyrki3 - 1):0]; 
assign Oztki3[0] = 1'b0; 
assign Oztki3[1] = (Zduki3[3:0] == 4'b0); 
assign Oztki3[2] = ((3 >= 2) ? (Deuki3[3:0] == 4'b0) : 1'b0); 
assign Oztki3[3] = ((3 >= 3) ? (Heuki3[3:0] == 4'b0) : 1'b0); 
assign Oztki3[4] = ((3 >= 4) ? (Leuki3[3:0] == 4'b0) : 1'b0); 
assign Oztki3[5] = ((3 >= 5) ? (Peuki3[3:0] == 4'b0) : 1'b0); 
assign Oztki3[6] = ((3 >= 6) ? (Teuki3[3:0] == 4'b0) : 1'b0); 
assign Oztki3[7] = ((3 >= 7) ? (Xeuki3[3:0] == 4'b0) : 1'b0); 
assign Oztki3[8] = ((3 >= 8) ? (Bfuki3[3:0] == 4'b0) : 1'b0); 
assign Oztki3[9] = ((3 >= 9) ? (Ffuki3[3:0] == 4'b0) : 1'b0); 
assign Oztki3[10] = ((3 >= 10) ? (Jfuki3[3:0] == 4'b0) : 1'b0); 
assign Oztki3[11] = ((3 >= 11) ? (Ofuki3[3:0] == 4'b0) : 1'b0); 
assign Oztki3[12] = ((3 >= 12) ? (Tfuki3[3:0] == 4'b0) : 1'b0); 
assign Oztki3[13] = ((3 >= 13) ? (Yfuki3[3:0] == 4'b0) : 1'b0); 
assign Oztki3[14] = ((3 >= 14) ? (Dguki3[3:0] == 4'b0) : 1'b0); 
assign Oztki3[15] = ((3 == 15) ? (Iguki3[3:0] == 4'b0) : 1'b0); 
assign H4ski3 = Oztki3[3:0]; 
assign D0uki3[3:0] = 4'hf; 
assign D0uki3[7:4] = (~Zduki3[3:0]); 
assign D0uki3[11:8] = (~Deuki3[3:0]); 
assign D0uki3[15:12] = (~Heuki3[3:0]); 
assign D0uki3[19:16] = (~Leuki3[3:0]); 
assign D0uki3[23:20] = (~Peuki3[3:0]); 
assign D0uki3[27:24] = (~Teuki3[3:0]); 
assign D0uki3[31:28] = (~Xeuki3[3:0]); 
assign D0uki3[35:32] = (~Bfuki3[3:0]); 
assign D0uki3[39:36] = (~Ffuki3[3:0]); 
assign D0uki3[43:40] = (~Jfuki3[3:0]); 
assign D0uki3[47:44] = (~Ofuki3[3:0]); 
assign D0uki3[51:48] = (~Tfuki3[3:0]); 
assign D0uki3[55:52] = (~Yfuki3[3:0]); 
assign D0uki3[59:56] = (~Dguki3[3:0]); 
assign D0uki3[63:60] = (~Iguki3[3:0]); 
assign S4ski3 = D0uki3[((4 * 4) - 1):0]; 
assign Yquki3 = Qjvki3; 
assign Nruki3 = ((3 >= 2) ? Dkvki3 : {32 {1'b0}}); 
assign Csuki3 = ((3 >= 3) ? Qkvki3 : {32 {1'b0}}); 
assign Rsuki3 = ((3 >= 4) ? Dlvki3 : {32 {1'b0}}); 
assign Gtuki3 = ((3 >= 5) ? Qlvki3 : {32 {1'b0}}); 
assign Vtuki3 = ((3 >= 6) ? Dmvki3 : {32 {1'b0}}); 
assign Kuuki3 = ((3 >= 7) ? Qmvki3 : {32 {1'b0}}); 
assign Zuuki3 = ((3 >= 8) ? Dnvki3 : {32 {1'b0}}); 
assign Ovuki3 = ((3 >= 9) ? Qnvki3 : {32 {1'b0}}); 
assign Dwuki3 = ((3 >= 10) ? Dovki3 : {32 {1'b0}}); 
assign Twuki3 = ((3 >= 11) ? Rovki3 : {32 {1'b0}}); 
assign Jxuki3 = ((3 >= 12) ? Fpvki3 : {32 {1'b0}}); 
assign Zxuki3 = ((3 >= 13) ? Tpvki3 : {32 {1'b0}}); 
assign Pyuki3 = ((3 >= 14) ? Hqvki3 : {32 {1'b0}}); 
assign Fzuki3 = ((3 >= 15) ? Vqvki3 : {32 {1'b0}}); 
assign F1tki3[(32 - 1):0] = Yquki3; 
assign F1tki3[((32 * 2) - 1):32] = Nruki3; 
assign F1tki3[((32 * 3) - 1):(32 * 2)] = Csuki3; 
assign F1tki3[((32 * 4) - 1):(32 * 3)] = Rsuki3; 
assign F1tki3[((32 * 5) - 1):(32 * 4)] = Gtuki3; 
assign F1tki3[((32 * 6) - 1):(32 * 5)] = Vtuki3; 
assign F1tki3[((32 * 7) - 1):(32 * 6)] = Kuuki3; 
assign F1tki3[((32 * 8) - 1):(32 * 7)] = Zuuki3; 
assign F1tki3[((32 * 9) - 1):(32 * 8)] = Ovuki3; 
assign F1tki3[((32 * 10) - 1):(32 * 9)] = Dwuki3; 
assign F1tki3[((32 * 11) - 1):(32 * 10)] = Twuki3; 
assign F1tki3[((32 * 12) - 1):(32 * 11)] = Jxuki3; 
assign F1tki3[((32 * 13) - 1):(32 * 12)] = Zxuki3; 
assign F1tki3[((32 * 14) - 1):(32 * 13)] = Pyuki3; 
assign F1tki3[((32 * 15) - 1):(32 * 14)] = Fzuki3; 
always @(posedge Yvrki3 or negedge Dwrki3) begin : H9wki3 
if (Dwrki3 == 1'b0) begin 
Qjuki3 <= 1'b0; 
end 
else 
begin 
if (Lwrki3 == 1'b1) begin 
Qjuki3 <= Keski3; 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : X9wki3 
if (Dwrki3 == 1'b0) begin 
Pkuki3 <= 32'b0; 
Zkuki3 <= 2'b0; 
Fjuki3 <= 1'b0; 
Kluki3 <= 3'b0; 
Dkuki3 <= 4'b0; 
end 
else 
begin 
if (Lwrki3 == 1'b1) begin 
Pkuki3 <= Peski3; 
Zkuki3 <= Swrki3; 
Fjuki3 <= Pfski3; 
Kluki3 <= Cfski3; 
Dkuki3 <= Qjski3; 
end 
end 
end 
always @(Peski3) begin : Fawki3 
Mquki3 = 1'b0; 
case (Peski3[9:0]) 
10'b0: 
Mquki3 = 1'b1; 
10'h004: 
if (3 > 1) begin 
Mquki3 = 1'b1; 
end 
10'h008: 
if (3 > 2) begin 
Mquki3 = 1'b1; 
end 
10'h00c: 
if (3 > 3) begin 
Mquki3 = 1'b1; 
end 
10'h010: 
if (3 > 4) begin 
Mquki3 = 1'b1; 
end 
10'h014: 
if (3 > 5) begin 
Mquki3 = 1'b1; 
end 
10'h018: 
if (3 > 6) begin 
Mquki3 = 1'b1; 
end 
10'h01c: 
if (3 > 7) begin 
Mquki3 = 1'b1; 
end 
10'h020: 
if (3 > 8) begin 
Mquki3 = 1'b1; 
end 
10'h024: 
if (3 > 9) begin 
Mquki3 = 1'b1; 
end 
10'h028: 
if (3 > 10) begin 
Mquki3 = 1'b1; 
end 
10'h02c: 
if (3 > 11) begin 
Mquki3 = 1'b1; 
end 
10'h030: 
if (3 > 12) begin 
Mquki3 = 1'b1; 
end 
10'h034: 
if (3 > 13) begin 
Mquki3 = 1'b1; 
end 
10'h038: 
if (3 > 14) begin 
Mquki3 = 1'b1; 
end 
10'h03c: 
if (1 == 1'b1) begin 
Mquki3 = 1'b1; 
end 
10'h040: 
if (1 == 1'b1) begin 
Mquki3 = 1'b1; 
end 
10'h044: 
if (1 == 1'b1) begin 
Mquki3 = 1'b1; 
end 
10'h048: 
Mquki3 = 1'b1; 
10'h04c: 
if (0 == 1'b1) begin 
Mquki3 = 1'b1; 
end 
10'h050: 
if (0 == 1'b1) begin 
Mquki3 = 1'b1; 
end 
10'h054: 
if (0 == 1'b1) begin 
Mquki3 = 1'b1; 
end 
10'h058: 
if ((0 == 1'b1) && (3 > 1)) begin 
Mquki3 = 1'b1; 
end 
10'h05c: 
if ((0 == 1'b1) && (3 > 2)) begin 
Mquki3 = 1'b1; 
end 
10'h060: 
if ((0 == 1'b1) && (3 > 3)) begin 
Mquki3 = 1'b1; 
end 
10'h064: 
if ((0 == 1'b1) && (3 > 4)) begin 
Mquki3 = 1'b1; 
end 
10'h068: 
if ((0 == 1'b1) && (3 > 5)) begin 
Mquki3 = 1'b1; 
end 
10'h06c: 
if ((0 == 1'b1) && (3 > 6)) begin 
Mquki3 = 1'b1; 
end 
10'h070: 
if ((0 == 1'b1) && (3 > 7)) begin 
Mquki3 = 1'b1; 
end 
10'h074: 
if ((0 == 1'b1) && (3 > 8)) begin 
Mquki3 = 1'b1; 
end 
10'h078: 
if ((0 == 1'b1) && (3 > 9)) begin 
Mquki3 = 1'b1; 
end 
10'h07c: 
if ((0 == 1'b1) && (3 > 10)) begin 
Mquki3 = 1'b1; 
end 
10'h080: 
if ((0 == 1'b1) && (3 > 11)) begin 
Mquki3 = 1'b1; 
end 
10'h084: 
if ((0 == 1'b1) && (3 > 12)) begin 
Mquki3 = 1'b1; 
end 
10'h088: 
if ((0 == 1'b1) && (3 > 13)) begin 
Mquki3 = 1'b1; 
end 
10'h08c: 
if ((0 == 1'b1) && (3 > 14)) begin 
Mquki3 = 1'b1; 
end 
10'h090: 
Mquki3 = 1'b1; 
default: 
Mquki3 = 1'b0; 
endcase 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Wawki3 
if (Dwrki3 == 1'b0) begin 
Uiuki3 <= 2'b0; 
end 
else 
begin 
if ((Fouki3 == Nauki3) || (Louki3 == Nauki3)) begin 
Uiuki3 <= 2'b1; 
end 
else begin 
Uiuki3 <= 2'b0; 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Mbwki3 
if (Dwrki3 == 1'b0) begin 
Nhuki3 <= 1'b1; 
end 
else begin 
Nhuki3 <= Eiuki3; 
end 
end 
always @(Fouki3 or Louki3 or Peski3 or Uluki3) begin : Gcwki3 
if ((((Fouki3 == Eauki3) && (Louki3 == W9uki3)) && (Peski3[9:0] == Uluki3[9:0])) 
|| (Louki3 == Nauki3)) begin 
Eiuki3 = 1'b0; 
end 
else begin 
Eiuki3 = 1'b1; 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Bdwki3 
if (Dwrki3 == 1'b0) begin 
Xnuki3 <= O9uki3; 
end 
else begin 
Xnuki3 <= Louki3; 
end 
end 
always @(Fouki3 or Hstki3 or Pfski3 or Mquki3 or Cfski3) begin : Mdwki3 
case (Fouki3) 
O9uki3, Eauki3, W9uki3: 
if (Hstki3 == 1'b1) begin 
if ((Mquki3 == 1'b1) && (Cfski3 == 3'b010)) begin 
if (Pfski3 == 1'b1) begin 
Louki3 = Eauki3; 
end 
else begin 
Louki3 = W9uki3; 
end 
end 
else begin 
Louki3 = Nauki3; 
end 
end 
else begin 
Louki3 = O9uki3; 
end 
default: 
Louki3 = O9uki3; 
endcase 
end 
always @(Ifski3 or Uluki3 or Z7wki3) begin : Bewki3 
if (Z7wki3 == 1'b1) begin 
if (Xyrki3 == 32) begin 
Vouki3 = Ifski3[31:0]; 
end 
else if (Xyrki3 == 64) begin 
case (Uluki3[2:0]) 
3'h4: 
Vouki3 = Ifski3[63:32]; 
default: 
Vouki3 = Ifski3[31:0]; 
endcase 
end 
else if (Xyrki3 == 128) begin 
case (Uluki3[3:0]) 
4'h4: 
Vouki3 = Ifski3[63:32]; 
4'h8: 
Vouki3 = Ifski3[95:64]; 
4'hc: 
Vouki3 = Ifski3[127:96]; 
default: 
Vouki3 = Ifski3[31:0]; 
endcase 
end 
else begin 
case (Uluki3[4:0]) 
5'h04: 
Vouki3 = Ifski3[63:32]; 
5'h08: 
Vouki3 = Ifski3[95:64]; 
5'h0c: 
Vouki3 = Ifski3[127:96]; 
5'h10: 
Vouki3 = Ifski3[159:128]; 
5'h14: 
Vouki3 = Ifski3[191:160]; 
5'h18: 
Vouki3 = Ifski3[223:192]; 
5'h1c: 
Vouki3 = Ifski3[255:224]; 
default: 
Vouki3 = Ifski3[31:0]; 
endcase 
end 
end 
else if (Xyrki3 == 32) begin 
Vouki3[7:0] = Ifski3[31:24]; 
Vouki3[15:8] = Ifski3[23:16]; 
Vouki3[23:16] = Ifski3[15:8]; 
Vouki3[31:24] = Ifski3[7:0]; 
end 
else if (Xyrki3 == 64) begin 
case (Uluki3[2:0]) 
3'h4: begin 
Vouki3[7:0] = Ifski3[31:24]; 
Vouki3[15:8] = Ifski3[23:16]; 
Vouki3[23:16] = Ifski3[15:8]; 
Vouki3[31:24] = Ifski3[7:0]; 
end 
default: begin 
Vouki3[7:0] = Ifski3[63:56]; 
Vouki3[15:8] = Ifski3[55:48]; 
Vouki3[23:16] = Ifski3[47:40]; 
Vouki3[31:24] = Ifski3[39:32]; 
end 
endcase 
end 
else if (Xyrki3 == 128) begin 
case (Uluki3[3:0]) 
4'h4: begin 
Vouki3[7:0] = Ifski3[95:88]; 
Vouki3[15:8] = Ifski3[87:80]; 
Vouki3[23:16] = Ifski3[79:72]; 
Vouki3[31:24] = Ifski3[71:64]; 
end 
4'h8: begin 
Vouki3[7:0] = Ifski3[63:56]; 
Vouki3[15:8] = Ifski3[55:48]; 
Vouki3[23:16] = Ifski3[47:40]; 
Vouki3[31:24] = Ifski3[39:32]; 
end 
4'hc: begin 
Vouki3[7:0] = Ifski3[31:24]; 
Vouki3[15:8] = Ifski3[23:16]; 
Vouki3[23:16] = Ifski3[15:8]; 
Vouki3[31:24] = Ifski3[7:0]; 
end 
default: begin 
Vouki3[7:0] = Ifski3[127:120]; 
Vouki3[15:8] = Ifski3[119:112]; 
Vouki3[23:16] = Ifski3[111:104]; 
Vouki3[31:24] = Ifski3[103:96]; 
end 
endcase 
end 
else begin 
case (Uluki3[4:0]) 
5'h04: begin 
Vouki3[7:0] = Ifski3[223:216]; 
Vouki3[15:8] = Ifski3[215:208]; 
Vouki3[23:16] = Ifski3[207:200]; 
Vouki3[31:24] = Ifski3[199:192]; 
end 
5'h08: begin 
Vouki3[7:0] = Ifski3[191:184]; 
Vouki3[15:8] = Ifski3[183:176]; 
Vouki3[23:16] = Ifski3[175:168]; 
Vouki3[31:24] = Ifski3[167:160]; 
end 
5'h0c: begin 
Vouki3[7:0] = Ifski3[159:152]; 
Vouki3[15:8] = Ifski3[151:144]; 
Vouki3[23:16] = Ifski3[143:136]; 
Vouki3[31:24] = Ifski3[135:128]; 
end 
5'h10: begin 
Vouki3[7:0] = Ifski3[127:120]; 
Vouki3[15:8] = Ifski3[119:112]; 
Vouki3[23:16] = Ifski3[111:104]; 
Vouki3[31:24] = Ifski3[103:96]; 
end 
5'h14: begin 
Vouki3[7:0] = Ifski3[95:88]; 
Vouki3[15:8] = Ifski3[87:80]; 
Vouki3[23:16] = Ifski3[79:72]; 
Vouki3[31:24] = Ifski3[71:64]; 
end 
5'h18: begin 
Vouki3[7:0] = Ifski3[63:56]; 
Vouki3[15:8] = Ifski3[55:48]; 
Vouki3[23:16] = Ifski3[47:40]; 
Vouki3[31:24] = Ifski3[39:32]; 
end 
5'h1c: begin 
Vouki3[7:0] = Ifski3[31:24]; 
Vouki3[15:8] = Ifski3[23:16]; 
Vouki3[23:16] = Ifski3[15:8]; 
Vouki3[31:24] = Ifski3[7:0]; 
end 
default: begin 
Vouki3[7:0] = Ifski3[255:248]; 
Vouki3[15:8] = Ifski3[247:240]; 
Vouki3[23:16] = Ifski3[239:232]; 
Vouki3[31:24] = Ifski3[231:224]; 
end 
endcase 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Rewki3 
if (Dwrki3 == 1'b0) begin 
Wauki3 <= 4'b1; 
end 
else 
begin 
if (Rstki3 == 1'b1) begin 
if ((Nnuki3 == 4'b1) && (U0uki3 == 0)) begin 
Wauki3 <= Wauki3; 
end 
else 
begin 
Wauki3 <= U0uki3; 
end 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Bfwki3 
if (Dwrki3 == 1'b0) begin 
Bbuki3 <= 4'h2; 
end 
else 
begin 
if (Zstki3 == 1'b1) begin 
if ((Nnuki3 == 4'h2) && (E1uki3 == 0)) begin 
Bbuki3 <= Bbuki3; 
end 
else 
begin 
Bbuki3 <= E1uki3; 
end 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Lfwki3 
if (Dwrki3 == 1'b0) begin 
Gbuki3 <= 4'h3; 
end 
else 
begin 
if (Httki3 == 1'b1) begin 
if ((Nnuki3 == 4'h3) && (O1uki3 == 0)) begin 
Gbuki3 <= Gbuki3; 
end 
else 
begin 
Gbuki3 <= O1uki3; 
end 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Vfwki3 
if (Dwrki3 == 1'b0) begin 
Lbuki3 <= 4'h4; 
end 
else 
begin 
if (Pttki3 == 1'b1) begin 
if ((Nnuki3 == 4'h4) && (Y1uki3 == 0)) begin 
Lbuki3 <= Lbuki3; 
end 
else 
begin 
Lbuki3 <= Y1uki3; 
end 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Fgwki3 
if (Dwrki3 == 1'b0) begin 
Qbuki3 <= 4'h5; 
end 
else 
begin 
if (Xttki3 == 1'b1) begin 
if ((Nnuki3 == 4'h5) && (I2uki3 == 0)) begin 
Qbuki3 <= Qbuki3; 
end 
else 
begin 
Qbuki3 <= I2uki3; 
end 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Pgwki3 
if (Dwrki3 == 1'b0) begin 
Vbuki3 <= 4'h6; 
end 
else 
begin 
if (Futki3 == 1'b1) begin 
if ((Nnuki3 == 4'h6) && (S2uki3 == 0)) begin 
Vbuki3 <= Vbuki3; 
end 
else 
begin 
Vbuki3 <= S2uki3; 
end 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Zgwki3 
if (Dwrki3 == 1'b0) begin 
Acuki3 <= 4'h7; 
end 
else 
begin 
if (Nutki3 == 1'b1) begin 
if ((Nnuki3 == 4'h7) && (C3uki3 == 0)) begin 
Acuki3 <= Acuki3; 
end 
else 
begin 
Acuki3 <= C3uki3; 
end 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Jhwki3 
if (Dwrki3 == 1'b0) begin 
Fcuki3 <= 4'h8; 
end 
else 
begin 
if (Vutki3 == 1'b1) begin 
if ((Nnuki3 == 4'h8) && (M3uki3 == 0)) begin 
Fcuki3 <= Fcuki3; 
end 
else 
begin 
Fcuki3 <= M3uki3; 
end 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Thwki3 
if (Dwrki3 == 1'b0) begin 
Kcuki3 <= 4'h9; 
end 
else 
begin 
if (Dvtki3 == 1'b1) begin 
if ((Nnuki3 == 4'h9) && (W3uki3 == 0)) begin 
Kcuki3 <= Kcuki3; 
end 
else 
begin 
Kcuki3 <= W3uki3; 
end 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Diwki3 
if (Dwrki3 == 1'b0) begin 
Pcuki3 <= 4'ha; 
end 
else 
begin 
if (Lvtki3 == 1'b1) begin 
if ((Nnuki3 == 4'ha) && (G4uki3 == 0)) begin 
Pcuki3 <= Pcuki3; 
end 
else 
begin 
Pcuki3 <= G4uki3; 
end 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Oiwki3 
if (Dwrki3 == 1'b0) begin 
Vcuki3 <= 4'hb; 
end 
else 
begin 
if (Uvtki3 == 1'b1) begin 
if ((Nnuki3 == 4'hb) && (R4uki3 == 0)) begin 
Vcuki3 <= Vcuki3; 
end 
else 
begin 
Vcuki3 <= R4uki3; 
end 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Ziwki3 
if (Dwrki3 == 1'b0) begin 
Bduki3 <= 4'hc; 
end 
else 
begin 
if (Dwtki3 == 1'b1) begin 
if ((Nnuki3 == 4'hc) && (C5uki3 == 0)) begin 
Bduki3 <= Bduki3; 
end 
else 
begin 
Bduki3 <= C5uki3; 
end 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Kjwki3 
if (Dwrki3 == 1'b0) begin 
Hduki3 <= 4'hd; 
end 
else 
begin 
if (Mwtki3 == 1'b1) begin 
if ((Nnuki3 == 4'hd) && (N5uki3 == 0)) begin 
Hduki3 <= Hduki3; 
end 
else 
begin 
Hduki3 <= N5uki3; 
end 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Vjwki3 
if (Dwrki3 == 1'b0) begin 
Nduki3 <= 4'he; 
end 
else 
begin 
if (Vwtki3 == 1'b1) begin 
if ((Nnuki3 == 4'he) && (Y5uki3 == 0)) begin 
Nduki3 <= Nduki3; 
end 
else 
begin 
Nduki3 <= Y5uki3; 
end 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Gkwki3 
if (Dwrki3 == 1'b0) begin 
Tduki3 <= 4'hf; 
end 
else 
begin 
if (Extki3 == 1'b1) begin 
if ((Nnuki3 == 4'hf) && (J6uki3 == 0)) begin 
Tduki3 <= Tduki3; 
end 
else 
begin 
Tduki3 <= J6uki3; 
end 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Rkwki3 
if (Dwrki3 == 1'b0) begin 
Nguki3 <= 10'b0; 
end 
else 
begin 
if (Nxtki3 == 1'b1) begin 
Nguki3 <= E7uki3; 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Glwki3 
if (Dwrki3 == 1'b0) begin 
Xguki3 <= 1'b0; 
end 
else 
begin 
if (Aytki3 == 1'b1) begin 
Xguki3 <= C9uki3; 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Slwki3 
if (Dwrki3 == 1'b0) begin 
Ehuki3 <= 0; 
end 
else 
begin 
if (Kytki3 == 1'b1) begin 
if (T7uki3 > 3) begin 
Ehuki3 <= {4 {1'b0}}; 
end 
else 
begin 
Ehuki3 <= T7uki3; 
end 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Fmwki3 
if (Dwrki3 == 1'b0) begin 
Aquki3 <= 1'b0; 
end 
else 
begin 
if (Kyski3 == 1'b1) begin 
Aquki3 <= 1'b1; 
end 
else 
begin 
if (Zxski3 == 1'b1) begin 
Aquki3 <= 1'b0; 
end 
end 
end 
end 
always @(Peski3 or Hstki3 or Pfski3) begin : Smwki3 
if (((Hstki3 == 1'b1) && (Pfski3 == 1'b0)) && (Peski3[9:0] == 10'h044)) begin 
Zxski3 = 1'b1; 
end 
else begin 
Zxski3 = 1'b0; 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Inwki3 
if (Dwrki3 == 1'b0) begin 
Vzuki3 <= 1'b0; 
end 
else 
begin 
if (M0vki3 == 1'b1) begin 
Vzuki3 <= B0vki3; 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Tnwki3 
if (Dwrki3 == 1'b0) begin 
Fbvki3 <= 32'h0000ffff; 
end 
else 
begin 
if (Acvki3 == 1'b1) begin 
Fbvki3 <= Havki3; 
end 
end 
end 
always @(Vavki3) begin 
Obvki3 = 32'b0; 
Obvki3[(32 - 1):0] = Vavki3; 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Howki3 
if (Dwrki3 == 1'b0) begin 
Mcvki3 <= 32'h0000000f; 
end 
else 
begin 
if (K1wki3 == 1'b1) begin 
Mcvki3 <= Jrvki3; 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Yowki3 
if (Dwrki3 == 1'b0) begin 
Ycvki3 <= 32'h0000000f; 
end 
else 
begin 
if (V1wki3 == 1'b1) begin 
Ycvki3 <= Asvki3; 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Ppwki3 
if (Dwrki3 == 1'b0) begin 
Kdvki3 <= 32'h0000000f; 
end 
else 
begin 
if (G2wki3 == 1'b1) begin 
Kdvki3 <= Rsvki3; 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Gqwki3 
if (Dwrki3 == 1'b0) begin 
Wdvki3 <= 32'h0000000f; 
end 
else 
begin 
if (R2wki3 == 1'b1) begin 
Wdvki3 <= Itvki3; 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Xqwki3 
if (Dwrki3 == 1'b0) begin 
Ievki3 <= 32'h0000000f; 
end 
else 
begin 
if (C3wki3 == 1'b1) begin 
Ievki3 <= Ztvki3; 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Orwki3 
if (Dwrki3 == 1'b0) begin 
Uevki3 <= 32'h0000000f; 
end 
else 
begin 
if (N3wki3 == 1'b1) begin 
Uevki3 <= Quvki3; 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Fswki3 
if (Dwrki3 == 1'b0) begin 
Gfvki3 <= 32'h0000000f; 
end 
else 
begin 
if (Y3wki3 == 1'b1) begin 
Gfvki3 <= Hvvki3; 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Wswki3 
if (Dwrki3 == 1'b0) begin 
Sfvki3 <= 32'h0000000f; 
end 
else 
begin 
if (J4wki3 == 1'b1) begin 
Sfvki3 <= Yvvki3; 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Ntwki3 
if (Dwrki3 == 1'b0) begin 
Egvki3 <= 32'h0000000f; 
end 
else 
begin 
if (U4wki3 == 1'b1) begin 
Egvki3 <= Pwvki3; 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Euwki3 
if (Dwrki3 == 1'b0) begin 
Qgvki3 <= 32'h0000000f; 
end 
else 
begin 
if (F5wki3 == 1'b1) begin 
Qgvki3 <= Gxvki3; 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Wuwki3 
if (Dwrki3 == 1'b0) begin 
Dhvki3 <= 32'h0000000f; 
end 
else 
begin 
if (R5wki3 == 1'b1) begin 
Dhvki3 <= Yxvki3; 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Ovwki3 
if (Dwrki3 == 1'b0) begin 
Qhvki3 <= 32'h0000000f; 
end 
else 
begin 
if (D6wki3 == 1'b1) begin 
Qhvki3 <= Qyvki3; 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Gwwki3 
if (Dwrki3 == 1'b0) begin 
Divki3 <= 32'h0000000f; 
end 
else 
begin 
if (P6wki3 == 1'b1) begin 
Divki3 <= Izvki3; 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Ywwki3 
if (Dwrki3 == 1'b0) begin 
Qivki3 <= 32'h0000000f; 
end 
else 
begin 
if (B7wki3 == 1'b1) begin 
Qivki3 <= A0wki3; 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Qxwki3 
if (Dwrki3 == 1'b0) begin 
Djvki3 <= 32'h0000000f; 
end 
else 
begin 
if (N7wki3 == 1'b1) begin 
Djvki3 <= S0wki3; 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Iywki3 
if (Dwrki3 == 1'b0) begin 
Opuki3 <= 32'b0; 
end 
else 
begin 
if ((Fouki3 == Nauki3) || (Louki3 == Nauki3)) begin 
Opuki3 <= 32'b0; 
end 
else 
begin 
if ((((Hstki3 == 1'b1) && (Pfski3 == 1'b0)) && (Eiuki3 == 1'b1)) || (((Q8uki3 == 
1'b1) && (Tmuki3 == 1'b0)) && (Iiski3 == 1'b0))) begin 
case (U6uki3) 
10'b0: 
Opuki3 <= {28'b0, Zduki3}; 
10'h004: 
Opuki3 <= {28'b0, Deuki3}; 
10'h008: 
Opuki3 <= {28'b0, Heuki3}; 
10'h00c: 
Opuki3 <= {28'b0, Leuki3}; 
10'h010: 
Opuki3 <= {28'b0, Peuki3}; 
10'h014: 
Opuki3 <= {28'b0, Teuki3}; 
10'h018: 
Opuki3 <= {28'b0, Xeuki3}; 
10'h01c: 
Opuki3 <= {28'b0, Bfuki3}; 
10'h020: 
Opuki3 <= {28'b0, Ffuki3}; 
10'h024: 
Opuki3 <= {28'b0, Jfuki3}; 
10'h028: 
Opuki3 <= {28'b0, Ofuki3}; 
10'h02c: 
Opuki3 <= {28'b0, Tfuki3}; 
10'h030: 
Opuki3 <= {28'b0, Yfuki3}; 
10'h034: 
Opuki3 <= {28'b0, Dguki3}; 
10'h038: 
Opuki3 <= {28'b0, Iguki3}; 
10'h03c: 
Opuki3 <= {22'b0, Stski3}; 
10'h040: 
Opuki3 <= {31'b0, Txski3}; 
10'h044: 
Opuki3 <= {31'b0, Iquki3}; 
10'h048: 
Opuki3 <= {24'b0, Buski3}; 
10'h04c: 
Opuki3 <= {31'b0, R1tki3}; 
10'h050: 
Opuki3 <= Obvki3; 
10'h054: 
Opuki3 <= V0vki3; 
10'h058: 
Opuki3 <= L1vki3; 
10'h05c: 
Opuki3 <= B2vki3; 
10'h060: 
Opuki3 <= R2vki3; 
10'h064: 
Opuki3 <= H3vki3; 
10'h068: 
Opuki3 <= X3vki3; 
10'h06c: 
Opuki3 <= N4vki3; 
10'h070: 
Opuki3 <= D5vki3; 
10'h074: 
Opuki3 <= T5vki3; 
10'h078: 
Opuki3 <= J6vki3; 
10'h07c: 
Opuki3 <= A7vki3; 
10'h080: 
Opuki3 <= R7vki3; 
10'h084: 
Opuki3 <= I8vki3; 
10'h088: 
Opuki3 <= Z8vki3; 
10'h08c: 
Opuki3 <= Q9vki3; 
10'h090: 
Opuki3 <= R8wki3; 
endcase 
end 
end 
end 
end 
always @(Opuki3) begin : Zywki3 
Gpuki3 = 32'b0; 
if (1 == 1) begin 
Gpuki3[31:0] = Opuki3[31:0]; 
end 
end 
always @(Yquki3) begin : Mzwki3 
V0vki3 = 32'b0; 
V0vki3[(32 - 1):0] = Yquki3; 
end 
always @(Nruki3) begin : H0xki3 
L1vki3 = 32'b0; 
L1vki3[(32 - 1):0] = Nruki3; 
end 
always @(Csuki3) begin : C1xki3 
B2vki3 = 32'b0; 
B2vki3[(32 - 1):0] = Csuki3; 
end 
always @(Rsuki3) begin : X1xki3 
R2vki3 = 32'b0; 
R2vki3[(32 - 1):0] = Rsuki3; 
end 
always @(Gtuki3) begin : S2xki3 
H3vki3 = 32'b0; 
H3vki3[(32 - 1):0] = Gtuki3; 
end 
always @(Vtuki3) begin : N3xki3 
X3vki3 = 32'b0; 
X3vki3[(32 - 1):0] = Vtuki3; 
end 
always @(Kuuki3) begin : I4xki3 
N4vki3 = 32'b0; 
N4vki3[(32 - 1):0] = Kuuki3; 
end 
always @(Zuuki3) begin : D5xki3 
D5vki3 = 32'b0; 
D5vki3[(32 - 1):0] = Zuuki3; 
end 
always @(Ovuki3) begin : Y5xki3 
T5vki3 = 32'b0; 
T5vki3[(32 - 1):0] = Ovuki3; 
end 
always @(Dwuki3) begin : T6xki3 
J6vki3 = 32'b0; 
J6vki3[(32 - 1):0] = Dwuki3; 
end 
always @(Twuki3) begin : P7xki3 
A7vki3 = 32'b0; 
A7vki3[(32 - 1):0] = Twuki3; 
end 
always @(Jxuki3) begin : L8xki3 
R7vki3 = 32'b0; 
R7vki3[(32 - 1):0] = Jxuki3; 
end 
always @(Zxuki3) begin : H9xki3 
I8vki3 = 32'b0; 
I8vki3[(32 - 1):0] = Zxuki3; 
end 
always @(Pyuki3) begin : Daxki3 
Z8vki3 = 32'b0; 
Z8vki3[(32 - 1):0] = Pyuki3; 
end 
always @(Fzuki3) begin : Zaxki3 
Q9vki3 = 32'b0; 
Q9vki3[(32 - 1):0] = Fzuki3; 
end 
endmodule 
module C9tki3(R1tki3, Tuski3, Ivski3, Ewski3, Vwski3, Zuski3, Lwski3); 
input R1tki3; 
input [3:0] Tuski3; 
input [3:0] Ivski3; 
input Ewski3; 
input Vwski3; 
output [3:0] Zuski3; 
output Lwski3; 
reg [3:0] Zuski3; 
reg Lwski3; 
always @(R1tki3 or Vwski3 or Ivski3 or Tuski3) begin 
Zuski3 = Tuski3; 
if (0 == 1) begin 
if ((R1tki3 == 1'b1) && (Vwski3 == 1'b0)) begin 
Zuski3 = Ivski3; 
end 
end 
end 
always @(R1tki3 or Vwski3 or Ewski3) begin 
Lwski3 = Ewski3; 
if (0 == 1) begin 
if (R1tki3 == 1'b1) begin 
Lwski3 = (Ewski3 && Vwski3); 
end 
end 
end 
endmodule 
module Vbxki3(Peski3, Hcxki3, Keski3); 
parameter Jsski3 = 32; 
`define Q5lkc `R1_N_SA_1
parameter Pcxki3 = `Q5lkc; 
`define T6lkc `R1_N_EA_1
parameter Zcxki3 = `T6lkc; 
`define K8lkc `R1_N_SA_2
parameter Jdxki3 = `K8lkc; 
`define E2lkc `R1_N_EA_2
parameter Tdxki3 = `E2lkc; 
input [(Jsski3 - 1):0] Peski3; 
input Hcxki3; 
output [(4 - 1):0] Keski3; 
wire [15:0] Dexki3; 
wire [15:0] Nexki3; 
wire [2:0] Afxki3; 
reg Zwrki3; 
integer P9ski3; 
`define N5lkc `R1_N_SA_0
assign Dexki3[0] = ((1 == 1) ? ((Peski3 >= `N5lkc) && (Peski3 <=  
`define R7lkc `R1_N_EA_0
`R7lkc)) : 1'b0); 
assign Dexki3[1] = ((((((((((Peski3 >= Pcxki3) && (Peski3 <= Zcxki3)) || ((( 
Peski3 >= 32'h03000000) && (Peski3 <= 32'h0300ffff)) && (0 >= 3'b1))) || ((( 
Peski3 >= 32'h04000000) && (Peski3 <= 32'h0400ffff)) && (0 >= 3'b010))) || ((( 
Peski3 >= 32'h05000000) && (Peski3 <= 32'h0500ffff)) && (0 >= 3'b011))) || ((( 
Peski3 >= 32'h06000000) && (Peski3 <= 32'h0600ffff)) && (0 >= 3'h4))) || ((( 
Peski3 >= 32'h07000000) && (Peski3 <= 32'h0700ffff)) && (0 >= 3'b101))) || ((( 
Peski3 >= 32'h08000000) && (Peski3 <= 32'h0800ffff)) && (0 >= 3'b110))) || ((( 
Peski3 >= 32'h09000000) && (Peski3 <= 32'h0900ffff)) && (0 == 3'b111))) && (1 != 
2'b10)); 
assign Dexki3[2] = ((((Peski3 >= Jdxki3) && (Peski3 <= Tdxki3)) || (((Peski3 >=  
`define O2lkc `R2_N_SA_2
`define W2lkc `R2_N_EA_2
`O2lkc) && (Peski3 <= `W2lkc)) && (0 == 1'b1))) && (1 != 2'b10)); 
assign Dexki3[3] = ((((Peski3 >= 32'h0c000000) && (Peski3 <= 32'h0c00ffff)) || ( 
((Peski3 >= 32'h0d000000) && (Peski3 <= 32'h0d00ffff)) && (0 == 1'b1))) && (1 != 
2'b10)); 
assign Dexki3[4] = ((((Peski3 >= 32'h0e000000) && (Peski3 <= 32'h0e00ffff)) || ( 
((Peski3 >= 32'h0f000000) && (Peski3 <= 32'h0f00ffff)) && (0 == 1'b1))) && (1 != 
2'b10)); 
assign Dexki3[5] = ((((Peski3 >= 32'h10000000) && (Peski3 <= 32'h1000ffff)) || ( 
((Peski3 >= 32'h11000000) && (Peski3 <= 32'h1100ffff)) && (0 == 1'b1))) && (1 != 
2'b10)); 
assign Dexki3[6] = ((((Peski3 >= 32'h12000000) && (Peski3 <= 32'h1200ffff)) || ( 
((Peski3 >= 32'h13000000) && (Peski3 <= 32'h1300ffff)) && (0 == 1'b1))) && (1 != 
2'b10)); 
assign Dexki3[7] = ((((Peski3 >= 32'h14000000) && (Peski3 <= 32'h1400ffff)) || ( 
((Peski3 >= 32'h15000000) && (Peski3 <= 32'h1500ffff)) && (0 == 1'b1))) && (1 != 
2'b10)); 
assign Dexki3[8] = ((((Peski3 >= 32'h16000000) && (Peski3 <= 32'h1600ffff)) || ( 
((Peski3 >= 32'h17000000) && (Peski3 <= 32'h1700ffff)) && (0 == 1'b1))) && (1 != 
2'b10)); 
assign Dexki3[9] = ((((Peski3 >= 32'h18000000) && (Peski3 <= 32'h1800ffff)) || ( 
((Peski3 >= 32'h19000000) && (Peski3 <= 32'h1900ffff)) && (0 == 1'b1))) && (1 != 
2'b10)); 
assign Dexki3[10] = ((((Peski3 >= 32'h1a000000) && (Peski3 <= 32'h1a00ffff)) ||  
(((Peski3 >= 32'h1b000000) && (Peski3 <= 32'h1b00ffff)) && (0 == 1'b1))) && (1  
!= 2'b10)); 
assign Dexki3[11] = ((((Peski3 >= 32'h1c000000) && (Peski3 <= 32'h1c00ffff)) ||  
(((Peski3 >= 32'h1d000000) && (Peski3 <= 32'h1d00ffff)) && (0 == 1'b1))) && (1  
!= 2'b10)); 
assign Dexki3[12] = ((((Peski3 >= 32'h1e000000) && (Peski3 <= 32'h1e00ffff)) ||  
(((Peski3 >= 32'h1f000000) && (Peski3 <= 32'h1f00ffff)) && (0 == 1'b1))) && (1  
!= 2'b10)); 
assign Dexki3[13] = ((((Peski3 >= 32'h20000000) && (Peski3 <= 32'h2000ffff)) ||  
(((Peski3 >= 32'h21000000) && (Peski3 <= 32'h2100ffff)) && (0 == 1'b1))) && (1  
!= 2'b10)); 
assign Dexki3[14] = ((((Peski3 >= 32'h22000000) && (Peski3 <= 32'h2200ffff)) ||  
(((Peski3 >= 32'h23000000) && (Peski3 <= 32'h2300ffff)) && (0 == 1'b1))) && (1  
!= 2'b10)); 
assign Dexki3[15] = ((((Peski3 >= 32'h24000000) && (Peski3 <= 32'h2400ffff)) ||  
(((Peski3 >= 32'h25000000) && (Peski3 <= 32'h2500ffff)) && (0 == 1'b1))) && (1  
!= 2'b10)); 
assign Nexki3[0] = ((1 == 1) ? ((Peski3 >= 32'h26000000) && (Peski3 <=  
32'h260003ff)) : 1'b0); 
assign Nexki3[1] = ((((((((((Peski3 >= 32'h27000000) && (Peski3 <= 32'h2700ffff) 
) || (((Peski3 >= 32'h28000000) && (Peski3 <= 32'h2800ffff)) && (0 >= 3'b1))) || 
(((Peski3 >= 32'h29000000) && (Peski3 <= 32'h2900ffff)) && (0 >= 3'b010))) || (( 
(Peski3 >= 32'h2a000000) && (Peski3 <= 32'h2a00ffff)) && (0 >= 3'b011))) || ((( 
Peski3 >= 32'h2b000000) && (Peski3 <= 32'h2b00ffff)) && (0 >= 3'h4))) || ((( 
Peski3 >= 32'h2c000000) && (Peski3 <= 32'h2c00ffff)) && (0 >= 3'b101))) || ((( 
Peski3 >= 32'h2d000000) && (Peski3 <= 32'h2d00ffff)) && (0 >= 3'b110))) || ((( 
Peski3 >= 32'h2e000000) && (Peski3 <= 32'h2e00ffff)) && (0 == 3'b111))) && (1 != 
2'b1)); 
assign Nexki3[2] = ((((Peski3 >= 32'h2f000000) && (Peski3 <= 32'h2f00ffff)) || ( 
((Peski3 >= 32'h30000000) && (Peski3 <= 32'h3000ffff)) && (0 == 1'b1))) && (1 != 
2'b1)); 
assign Nexki3[3] = ((((Peski3 >= 32'h31000000) && (Peski3 <= 32'h3100ffff)) || ( 
((Peski3 >= 32'h32000000) && (Peski3 <= 32'h3200ffff)) && (0 == 1'b1))) && (1 != 
2'b1)); 
assign Nexki3[4] = ((((Peski3 >= 32'h33000000) && (Peski3 <= 32'h3300ffff)) || ( 
((Peski3 >= 32'h34000000) && (Peski3 <= 32'h3400ffff)) && (0 == 1'b1))) && (1 != 
2'b1)); 
assign Nexki3[5] = ((((Peski3 >= 32'h35000000) && (Peski3 <= 32'h3500ffff)) || ( 
((Peski3 >= 32'h36000000) && (Peski3 <= 32'h3600ffff)) && (0 == 1'b1))) && (1 != 
2'b1)); 
assign Nexki3[6] = ((((Peski3 >= 32'h37000000) && (Peski3 <= 32'h3700ffff)) || ( 
((Peski3 >= 32'h38000000) && (Peski3 <= 32'h3800ffff)) && (0 == 1'b1))) && (1 != 
2'b1)); 
assign Nexki3[7] = ((((Peski3 >= 32'h39000000) && (Peski3 <= 32'h3900ffff)) || ( 
((Peski3 >= 32'h3a000000) && (Peski3 <= 32'h3a00ffff)) && (0 == 1'b1))) && (1 != 
2'b1)); 
assign Nexki3[8] = ((((Peski3 >= 32'h3b000000) && (Peski3 <= 32'h3b00ffff)) || ( 
((Peski3 >= 32'h3c000000) && (Peski3 <= 32'h3c00ffff)) && (0 == 1'b1))) && (1 != 
2'b1)); 
assign Nexki3[9] = ((((Peski3 >= 32'h3d000000) && (Peski3 <= 32'h3d00ffff)) || ( 
((Peski3 >= 32'h3e000000) && (Peski3 <= 32'h3e00ffff)) && (0 == 1'b1))) && (1 != 
2'b1)); 
assign Nexki3[10] = ((((Peski3 >= 32'h3f000000) && (Peski3 <= 32'h3f00ffff)) ||  
(((Peski3 >= 32'h40000000) && (Peski3 <= 32'h4000ffff)) && (0 == 1'b1))) && (1  
!= 2'b1)); 
assign Nexki3[11] = ((((Peski3 >= 32'h41000000) && (Peski3 <= 32'h4100ffff)) ||  
(((Peski3 >= 32'h42000000) && (Peski3 <= 32'h4200ffff)) && (0 == 1'b1))) && (1  
!= 2'b1)); 
assign Nexki3[12] = ((((Peski3 >= 32'h43000000) && (Peski3 <= 32'h4300ffff)) ||  
(((Peski3 >= 32'h44000000) && (Peski3 <= 32'h4400ffff)) && (0 == 1'b1))) && (1  
!= 2'b1)); 
assign Nexki3[13] = ((((Peski3 >= 32'h45000000) && (Peski3 <= 32'h4500ffff)) ||  
(((Peski3 >= 32'h46000000) && (Peski3 <= 32'h4600ffff)) && (0 == 1'b1))) && (1  
!= 2'b1)); 
assign Nexki3[14] = ((((Peski3 >= 32'h47000000) && (Peski3 <= 32'h4700ffff)) ||  
(((Peski3 >= 32'h48000000) && (Peski3 <= 32'h4800ffff)) && (0 == 1'b1))) && (1  
!= 2'b1)); 
assign Nexki3[15] = ((((Peski3 >= 32'h49000000) && (Peski3 <= 32'h4900ffff)) ||  
(((Peski3 >= 32'h4a000000) && (Peski3 <= 32'h4a00ffff)) && (0 == 1'b1))) && (1  
!= 2'b1)); 
assign Afxki3 = (Hcxki3 ? Dexki3[2:0] : Nexki3[2:0]); 
assign Keski3[2:0] = Afxki3; 
assign Keski3[(2 + 1)] = Zwrki3; 
always @(Afxki3) begin : Jfxki3 
Zwrki3 = 1'b1; 
for (P9ski3 = 0; (P9ski3 <= 2); P9ski3 = (P9ski3 + 1)) begin 
if (Afxki3[P9ski3] == 1'b1) begin 
Zwrki3 = 1'b0; 
end 
end 
end 
endmodule 
module K5tki3(Yvrki3, Dwrki3, Zdski3, Veski3, Lwrki3, D3ski3, U5ski3, Swrki3,  
Wfski3, Buski3, Sgski3, Zuski3, Lwski3, B6ski3, Kyski3, Ggski3, O2tki3, S0tki3,  
F5ski3, K5ski3, Nhski3, Yjski3, Qjski3, Syski3, Q5ski3); 
parameter Yfxki3 = 2'b0; 
parameter Agxki3 = 2'b1; 
parameter Cgxki3 = 2'b10; 
parameter Fgxki3 = 2'b11; 
input Yvrki3; 
input Dwrki3; 
input Zdski3; 
input [(3 - 1):0] Veski3; 
input Lwrki3; 
input [(2 - 1):0] D3ski3; 
input [(16 - 1):0] U5ski3; 
input [(2 - 1):0] Swrki3; 
input [3:0] Wfski3; 
input [3:0] Ggski3; 
input [(4 - 1):0] Buski3; 
input Sgski3; 
input [3:0] Zuski3; 
input Lwski3; 
input [3:0] B6ski3; 
input Kyski3; 
output O2tki3; 
output [3:0] S0tki3; 
output F5ski3; 
output K5ski3; 
output [3:0] Nhski3; 
output Yjski3; 
output [(4 - 1):0] Qjski3; 
output Syski3; 
output Q5ski3; 
reg K5ski3; 
reg [3:0] Nhski3; 
reg [(4 - 1):0] Qjski3; 
reg Syski3; 
reg [15:0] Hgxki3; 
reg Ygxki3; 
reg Jhxki3; 
reg Thxki3; 
reg [1:0] Aixki3; 
reg [1:0] Iixki3; 
reg [(4 - 1):0] Nnuki3; 
reg [(4 - 1):0] Uixki3; 
reg Gjxki3; 
reg [3:0] Mjxki3; 
reg [3:0] Tjxki3; 
reg [3:0] Bkxki3; 
reg [3:0] Ekxki3; 
reg Ikxki3; 
reg [3:0] Pkxki3; 
reg [15:0] Flxki3; 
wire [3:0] Rlxki3; 
wire Cmxki3; 
wire Imxki3; 
wire Qmxki3; 
wire Vmxki3; 
wire Dnxki3; 
wire Knxki3; 
wire Pnxki3; 
wire Tnxki3; 
wire Goxki3; 
wire Koxki3; 
wire Soxki3; 
wire Zoxki3; 
integer P9ski3; 
integer R9ski3; 
integer Gpxki3; 
integer Ipxki3; 
assign Tnxki3 = (((Kyski3 == 1'b1) && (F5ski3 == 1'b0)) && (O2tki3 == 1'b0)); 
assign Pnxki3 = ((Lwrki3 == 1'b1) && ((Swrki3 == 2'b11) || (Swrki3 == 2'b10))); 
assign S0tki3 = Hgxki3[3:0]; 
assign O2tki3 = ((((Nhski3[0] == 1'b0) && (Pkxki3 != Nhski3)) && (Lwrki3 == 1'b1 
)) && (Zdski3 == 1'b0)); 
assign Koxki3 = (((Veski3 > 3'b1) && (Swrki3 == 2'b11)) && (D3ski3 == 2'b0)); 
assign Q5ski3 = ((Uixki3 == Nnuki3) && (Aixki3 == Fgxki3)); 
assign Qmxki3 = (Iixki3 != Yfxki3); 
assign Cmxki3 = ((Mjxki3 == 4'b0) && (Koxki3 == 1'b0)); 
assign Imxki3 = ((Mjxki3 == 4'b1) && (Lwrki3 == 1'b1)); 
assign Dnxki3 = (((((Qmxki3 == 1'b1) && (D3ski3 == 2'b11)) && (Aixki3 != Yfxki3) 
) && (K5ski3 == 1'b0)) || ((Qmxki3 == 1'b0) && ((Swrki3 != 2'b1) || (Cmxki3 ==  
1'b1)))); 
assign Goxki3 = ((((D3ski3 == 2'b10) || (D3ski3 == 2'b11)) && (Iixki3 == Yfxki3) 
) && (Lwrki3 == 1'b0)); 
assign Vmxki3 = ((((((((Imxki3 == 1'b1) || (Cmxki3 == 1'b1)) && (Dnxki3 == 1'b1) 
) && (O2tki3 == 1'b0)) || (((Aixki3 == Yfxki3) && (Iixki3 == Yfxki3)) && (Zdski3 
== 1'b1))) || (Goxki3 == 1'b1)) || (Aixki3 == Fgxki3)) || (Zoxki3 == 1'b1)); 
assign Rlxki3 = {{3 {1'b0}}, 1'b1}; 
assign Soxki3 = ((Sgski3 == 1'b1) && (Swrki3 == 2'b0)); 
assign Zoxki3 = ((1 == 1'b1) ? Soxki3 : Sgski3); 
assign Knxki3 = (((Lwrki3 == 1'b1) && (Ikxki3 == 1'b1)) || (Aixki3 == Cgxki3)); 
assign Yjski3 = (Aixki3 == Agxki3); 
assign F5ski3 = (Iixki3 != Yfxki3); 
always @(Wfski3 or Uixki3 or Jhxki3) begin : Kpxki3 
Ygxki3 = 1'b0; 
for (P9ski3 = 0; (P9ski3 <= 3); P9ski3 = (P9ski3 + 1)) begin 
Ygxki3 = ((((Wfski3[P9ski3] == 1'b1) && (Uixki3 == P9ski3)) && (Jhxki3 == 1'b1)) 
|| Ygxki3); 
end 
end 
always @(Lwrki3 or Aixki3) begin : Aqxki3 
if (Aixki3 == Fgxki3) begin 
Jhxki3 = 1'b0; 
end 
else 
begin 
Jhxki3 = Lwrki3; 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Pqxki3 
if (Dwrki3 == 1'b0) begin 
Thxki3 <= 1'b0; 
end 
else 
begin 
if (Jhxki3 == 1'b1) begin 
Thxki3 <= Ygxki3; 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Brxki3 
if (Dwrki3 == 1'b0) begin 
Gjxki3 <= 1'b0; 
end 
else 
begin 
if (Aixki3 == Fgxki3) begin 
Gjxki3 <= 1'b1; 
end 
else begin 
Gjxki3 <= 1'b0; 
end 
end 
end 
always @(D3ski3 or Swrki3 or Veski3 or Bkxki3 or Tnxki3 or Lwrki3 or Zdski3)  
begin : Mrxki3 
if (((((((((Tnxki3 == 1'b1) || ((D3ski3 == 2'b11) && (Lwrki3 == 1'b0))) || (( 
D3ski3 == 2'b10) && (Lwrki3 == 1'b0))) || ((D3ski3 == 2'b11) && (Swrki3 == 2'b0) 
)) || ((D3ski3 == 2'b10) && (Swrki3 == 2'b0))) || (Swrki3 == 2'b0)) || (Zdski3  
== 1'b1)) || ((Veski3 == 3'b1) && (0 == 0))) || (Veski3 == 3'b0)) begin 
Mjxki3 = 4'b0; 
end 
else 
begin 
if (((Veski3 == 3'b111) || (Veski3 == 3'b110)) && (Swrki3 == 2'b10)) begin 
Mjxki3 = 4'hf; 
end 
else 
begin 
if (((Veski3 == 3'b101) || (Veski3 == 3'h4)) && (Swrki3 == 2'b10)) begin 
Mjxki3 = 4'h7; 
end 
else 
begin 
if (((Veski3 == 3'b011) || (Veski3 == 3'b010)) && (Swrki3 == 2'b10)) begin 
Mjxki3 = 4'h3; 
end 
else 
begin 
if ((Veski3 == 3'b1) && (0 == 1)) begin 
Mjxki3 = 4'hf; 
end 
else 
begin 
if (Bkxki3 == 4'b0) begin 
Mjxki3 = 4'b0; 
end 
else 
begin 
Mjxki3 = (Bkxki3 - 4'b1); 
end 
end 
end 
end 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Yrxki3 
if (Dwrki3 == 1'b0) begin 
Bkxki3 <= 4'b0; 
end 
else 
begin 
if (Pnxki3 == 1'b1) begin 
Bkxki3 <= Mjxki3; 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Gsxki3 
if (Dwrki3 == 1'b0) begin 
Pkxki3 <= {4 {1'b1}}; 
end 
else 
begin 
Pkxki3 <= Nhski3; 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Usxki3 
if (Dwrki3 == 1'b0) begin 
Ekxki3 <= 4'b0; 
end 
else 
begin 
if (Pnxki3 == 1'b1) begin 
Ekxki3 <= Tjxki3; 
end 
end 
end 
always @(Veski3 or Swrki3 or Ekxki3) begin : Dtxki3 
if (Veski3 > 3'b1) begin 
case (Swrki3) 
2'b10: 
case (Veski3[2:1]) 
1: 
Tjxki3 = 4'h3; 
2: 
Tjxki3 = 4'h7; 
default: 
Tjxki3 = 4'hf; 
endcase 
2'b11: 
Tjxki3 = (Ekxki3 - 4'b1); 
2'b0: 
Tjxki3 = 4'b0; 
default: 
Tjxki3 = Ekxki3; 
endcase 
end 
else 
begin 
Tjxki3 = 4'b0; 
end 
end 
always @(Tjxki3 or Ggski3 or Qjski3) begin : Qtxki3 
Hgxki3 = Ggski3; 
if (Tjxki3 > 4'b1) begin 
Hgxki3[Qjski3] = 1'b1; 
end 
end 
always @(B6ski3) begin : Euxki3 
Flxki3 <= 16'b0; 
Flxki3[3:0] <= B6ski3; 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Vuxki3 
if (Dwrki3 == 1'b0) begin 
Nhski3 <= {{3 {1'b0}}, 1'b1}; 
end 
else if (Vmxki3 == 1'b1) begin 
if (((((Qmxki3 == 1'b1) && (D3ski3 == 2'b11)) && (Lwrki3 == 1'b0)) || (Tnxki3 == 
1'b1)) || (Zoxki3 == 1'b1)) begin 
Nhski3 <= Rlxki3; 
end 
else 
begin 
if ((Aixki3 == Cgxki3) && (D3ski3 == 2'b10)) begin 
for (R9ski3 = 0; (R9ski3 <= 3); R9ski3 = (R9ski3 + 1)) begin 
Nhski3[R9ski3] <= (Nnuki3 == R9ski3[3:0]); 
end 
end 
else 
begin 
if (Lwski3 == 1'b1) begin 
if ((D3ski3 == 2'b10) && (Lwrki3 == 1'b0)) begin 
for (R9ski3 = 0; (R9ski3 <= 3); R9ski3 = (R9ski3 + 1)) begin 
Nhski3[R9ski3] <= (Nnuki3 == R9ski3[3:0]); 
end 
end 
else 
begin 
if (Flxki3[Buski3] == 1'b1) begin 
Nhski3 <= Rlxki3; 
end 
else 
begin 
for (R9ski3 = 0; (R9ski3 <= 3); R9ski3 = (R9ski3 + 1)) begin 
Nhski3[R9ski3] <= (Buski3 == R9ski3[3:0]); 
end 
end 
end 
end 
else 
begin 
Nhski3 <= Zuski3; 
end 
end 
end 
end 
else 
begin 
if (Tnxki3 == 1'b1) begin 
Nhski3 <= Rlxki3; 
end 
end 
end 
always @(Nhski3 or Buski3) begin : Lvxki3 
Uixki3 = Buski3; 
for (Gpxki3 = 0; (Gpxki3 <= 3); Gpxki3 = (Gpxki3 + 1)) begin 
if (Nhski3[Gpxki3] == 1'b1) begin 
Uixki3 = Gpxki3[3:0]; 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Cwxki3 
if (Dwrki3 == 1'b0) begin 
Qjski3 <= {4 {1'b0}}; 
end 
else 
begin 
if (Lwrki3 == 1'b1) begin 
Qjski3 <= Uixki3; 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Pwxki3 
if (Dwrki3 == 1'b0) begin 
Ikxki3 <= 1'b0; 
end 
else 
begin 
if (Lwrki3 == 1'b1) begin 
if (Aixki3 == Yfxki3) begin 
Ikxki3 <= 1'b1; 
end 
else 
begin 
Ikxki3 <= 1'b0; 
end 
end 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Bxxki3 
if (Dwrki3 == 1'b0) begin 
Nnuki3 <= {4 {1'b0}}; 
end 
else 
begin 
if (Knxki3 == 1'b1) begin 
Nnuki3 <= Qjski3; 
end 
end 
end 
always @(Swrki3 or Thxki3) begin : Qxxki3 
if (((Swrki3 == 2'b10) || (Swrki3 == 2'b0)) || (Thxki3 == 1'b1)) begin 
Syski3 = 1'b1; 
end 
else begin 
Syski3 = 1'b0; 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Dyxki3 
if (Dwrki3 == 1'b0) begin 
Aixki3 <= Yfxki3; 
end 
else begin 
Aixki3 <= Iixki3; 
end 
end 
always @(Aixki3 or Lwrki3 or Ygxki3 or Thxki3 or Swrki3 or Gjxki3 or D3ski3 or  
Uixki3 or Nnuki3 or K5ski3 or Qjski3) begin : Qyxki3 
case (Aixki3) 
Agxki3: 
if ((Lwrki3 == 1'b1) && (Swrki3 != 2'b1)) begin 
if ((Ygxki3 == 1'b1) || ((Thxki3 == 1'b1) && (Gjxki3 == 1'b1))) begin 
Iixki3 = Agxki3; 
end 
else begin 
Iixki3 = Cgxki3; 
end 
end 
else 
begin 
if ((D3ski3 == 2'b11) && (K5ski3 == 1'b0)) begin 
Iixki3 = Fgxki3; 
end 
else 
begin 
if (((K5ski3 == 1'b1) && (Qjski3 == Nnuki3)) && ((D3ski3 == 2'b10) || (D3ski3 == 
2'b11))) begin 
Iixki3 = Yfxki3; 
end 
else 
begin 
Iixki3 = Agxki3; 
end 
end 
end 
Cgxki3: 
if ((Lwrki3 == 1'b1) && (Swrki3 != 2'b1)) begin 
if ((Ygxki3 == 1'b1) || (D3ski3 == 2'b10)) begin 
Iixki3 = Agxki3; 
end 
else begin 
Iixki3 = Yfxki3; 
end 
end 
else 
begin 
if (D3ski3 == 2'b11) begin 
Iixki3 = Fgxki3; 
end 
else begin 
Iixki3 = Cgxki3; 
end 
end 
Fgxki3: 
if ((Lwrki3 == 1'b1) && (Uixki3 == Nnuki3)) begin 
Iixki3 = Agxki3; 
end 
else begin 
Iixki3 = Fgxki3; 
end 
default: 
if ((Lwrki3 == 1'b1) && (Ygxki3 == 1'b1)) begin 
Iixki3 = Agxki3; 
end 
else 
begin 
Iixki3 = Yfxki3; 
end 
endcase 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin 
if (Dwrki3 == 1'b0) begin 
K5ski3 <= 1'b0; 
end 
else 
begin 
if ((Aixki3 == Yfxki3) && (Iixki3 == Agxki3)) begin 
K5ski3 <= 1'b1; 
end 
else 
begin 
if (Lwrki3 == 1'b1) begin 
K5ski3 <= 1'b0; 
end 
end 
end 
end 
endmodule 
module Izxki3(Yvrki3, Dwrki3, Lwrki3, Qjski3, Sgski3, R1tki3, W1tki3, F1tki3,  
B6ski3, Ikski3, Vkski3, Ilski3, Vlski3, Imski3, Vmski3, Inski3, Unski3, Goski3,  
Soski3, Epski3, Qpski3, Cqski3, Oqski3, Arski3, Juski3, Yrski3); 
input Yvrki3; 
input Dwrki3; 
input Lwrki3; 
input Sgski3; 
input R1tki3; 
input [3:0] B6ski3; 
input [(4 - 1):0] Qjski3; 
input [(32 - 1):0] W1tki3; 
input [(480 - 1):0] F1tki3; 
output [(32 - 1):0] Ikski3; 
output [(32 - 1):0] Vkski3; 
output [(32 - 1):0] Ilski3; 
output [(32 - 1):0] Vlski3; 
output [(32 - 1):0] Imski3; 
output [(32 - 1):0] Vmski3; 
output [(32 - 1):0] Inski3; 
output [(32 - 1):0] Unski3; 
output [(32 - 1):0] Goski3; 
output [(32 - 1):0] Soski3; 
output [(32 - 1):0] Epski3; 
output [(32 - 1):0] Qpski3; 
output [(32 - 1):0] Cqski3; 
output [(32 - 1):0] Oqski3; 
output [(32 - 1):0] Arski3; 
output [3:0] Juski3; 
output Yrski3; 
reg [(32 - 1):0] Uzxki3; 
wire [15:0] E0yki3; 
wire [(32 - 1):0] M0yki3; 
wire [(32 - 1):0] A1yki3; 
wire [(32 - 1):0] O1yki3; 
wire [(32 - 1):0] C2yki3; 
wire [(32 - 1):0] Q2yki3; 
wire [(32 - 1):0] E3yki3; 
wire [(32 - 1):0] S3yki3; 
wire [(32 - 1):0] F4yki3; 
wire [(32 - 1):0] S4yki3; 
wire [(32 - 1):0] F5yki3; 
wire [(32 - 1):0] S5yki3; 
wire [(32 - 1):0] F6yki3; 
wire [(32 - 1):0] S6yki3; 
wire [(32 - 1):0] F7yki3; 
wire [(32 - 1):0] S7yki3; 
wire F8yki3; 
wire O8yki3; 
wire B9yki3; 
wire Q9yki3; 
wire Fayki3; 
wire Uayki3; 
wire Jbyki3; 
wire Ybyki3; 
wire Ncyki3; 
wire Cdyki3; 
wire Rdyki3; 
wire Geyki3; 
wire Weyki3; 
wire Mfyki3; 
wire Cgyki3; 
wire Sgyki3; 
wire Ihyki3; 
wire Yhyki3; 
wire Jiyki3; 
wire Uiyki3; 
wire Fjyki3; 
wire Qjyki3; 
wire Bkyki3; 
wire Mkyki3; 
wire Xkyki3; 
wire Ilyki3; 
wire Tlyki3; 
wire Fmyki3; 
wire Rmyki3; 
wire Dnyki3; 
wire Pnyki3; 
wire Boyki3; 
wire Noyki3; 
wire Zoyki3; 
wire Lpyki3; 
wire Xpyki3; 
wire Jqyki3; 
wire Vqyki3; 
wire Hryki3; 
wire Tryki3; 
wire Fsyki3; 
wire Rsyki3; 
wire Etyki3; 
wire Rtyki3; 
wire Euyki3; 
wire Ruyki3; 
wire Evyki3; 
wire Rvyki3; 
reg Cwyki3; 
wire Kwyki3; 
wire Uwyki3; 
wire Fxyki3; 
reg Oxyki3; 
assign Yrski3 = Rvyki3; 
assign Fxyki3 = ((Oxyki3 == 1'b0) && (R1tki3 == 1'b1)); 
assign Kwyki3 = ((Cwyki3 == 1'b1) && (Sgski3 == 1'b0)); 
assign Uwyki3 = ((1 == 0) ? 1'b0 : Kwyki3); 
assign Rvyki3 = (((Uzxki3 == {32 {1'b0}}) || (Kwyki3 == 1'b1)) || (Fxyki3 ==  
1'b1)); 
assign F8yki3 = ((0 == 1'b0) ? 1'b1 : Lwrki3); 
assign O8yki3 = (R1tki3 && F8yki3); 
assign B9yki3 = ((Qjski3 == 4'b1) && (O8yki3 == 1'b1)); 
assign Noyki3 = ((0 == 1) ? Yhyki3 : 1'b0); 
assign Arski3 = ((0 == 1) ? S7yki3 : {32 {1'b0}}); 
assign Q9yki3 = ((Qjski3 == 4'h2) && (O8yki3 == 1'b1)); 
assign Zoyki3 = (((0 == 1) && (3 > 1)) ? Jiyki3 : 1'b0); 
assign Oqski3 = (((0 == 1) && (3 > 1)) ? F7yki3 : {32 {1'b0}}); 
assign Fayki3 = ((Qjski3 == 4'h3) && (O8yki3 == 1'b1)); 
assign Lpyki3 = (((0 == 1) && (3 > 2)) ? Uiyki3 : 1'b0); 
assign Cqski3 = (((0 == 1) && (3 > 2)) ? S6yki3 : {32 {1'b0}}); 
assign Uayki3 = ((Qjski3 == 4'h4) && (O8yki3 == 1'b1)); 
assign Xpyki3 = (((0 == 1) && (3 > 3)) ? Fjyki3 : 1'b0); 
assign Qpski3 = (((0 == 1) && (3 > 3)) ? F6yki3 : {32 {1'b0}}); 
assign Jbyki3 = ((Qjski3 == 4'h5) && (O8yki3 == 1'b1)); 
assign Jqyki3 = (((0 == 1) && (3 > 4)) ? Qjyki3 : 1'b0); 
assign Epski3 = (((0 == 1) && (3 > 4)) ? S5yki3 : {32 {1'b0}}); 
assign Ybyki3 = ((Qjski3 == 4'h6) && (O8yki3 == 1'b1)); 
assign Vqyki3 = (((0 == 1) && (3 > 5)) ? Bkyki3 : 1'b0); 
assign Soski3 = (((0 == 1) && (3 > 5)) ? F5yki3 : {32 {1'b0}}); 
assign Ncyki3 = ((Qjski3 == 4'h7) && (O8yki3 == 1'b1)); 
assign Hryki3 = (((0 == 1) && (3 > 6)) ? Mkyki3 : 1'b0); 
assign Goski3 = (((0 == 1) && (3 > 6)) ? S4yki3 : {32 {1'b0}}); 
assign Cdyki3 = ((Qjski3 == 4'h8) && (O8yki3 == 1'b1)); 
assign Tryki3 = (((0 == 1) && (3 > 7)) ? Xkyki3 : 1'b0); 
assign Unski3 = (((0 == 1) && (3 > 7)) ? F4yki3 : {32 {1'b0}}); 
assign Rdyki3 = ((Qjski3 == 4'h9) && (O8yki3 == 1'b1)); 
assign Fsyki3 = (((0 == 1) && (3 > 8)) ? Ilyki3 : 1'b0); 
assign Inski3 = (((0 == 1) && (3 > 8)) ? S3yki3 : {32 {1'b0}}); 
assign Geyki3 = ((Qjski3 == 4'ha) && (O8yki3 == 1'b1)); 
assign Rsyki3 = (((0 == 1) && (3 > 9)) ? Tlyki3 : 1'b0); 
assign Vmski3 = (((0 == 1) && (3 > 9)) ? E3yki3 : {32 {1'b0}}); 
assign Weyki3 = ((Qjski3 == 4'hb) && (O8yki3 == 1'b1)); 
assign Etyki3 = (((0 == 1) && (3 > 10)) ? Fmyki3 : 1'b0); 
assign Imski3 = (((0 == 1) && (3 > 10)) ? Q2yki3 : {32 {1'b0}}); 
assign Mfyki3 = ((Qjski3 == 4'hc) && (O8yki3 == 1'b1)); 
assign Rtyki3 = (((0 == 1) && (3 > 11)) ? Rmyki3 : 1'b0); 
assign Vlski3 = (((0 == 1) && (3 > 11)) ? C2yki3 : {32 {1'b0}}); 
assign Cgyki3 = ((Qjski3 == 4'hd) && (O8yki3 == 1'b1)); 
assign Euyki3 = (((0 == 1) && (3 > 12)) ? Dnyki3 : 1'b0); 
assign Ilski3 = (((0 == 1) && (3 > 12)) ? O1yki3 : {32 {1'b0}}); 
assign Sgyki3 = ((Qjski3 == 4'he) && (O8yki3 == 1'b1)); 
assign Ruyki3 = (((0 == 1) && (3 > 13)) ? Pnyki3 : 1'b0); 
assign Vkski3 = (((0 == 1) && (3 > 13)) ? A1yki3 : {32 {1'b0}}); 
assign Ihyki3 = ((Qjski3 == 4'hf) && (O8yki3 == 1'b1)); 
assign Evyki3 = (((0 == 1) && (3 > 14)) ? Boyki3 : 1'b0); 
assign Ikski3 = (((0 == 1) && (3 > 14)) ? M0yki3 : {32 {1'b0}}); 
assign E0yki3 = {Evyki3, Ruyki3, Euyki3, Rtyki3, Etyki3, Rsyki3, Fsyki3, Tryki3, 
Hryki3, Vqyki3, Jqyki3, Xpyki3, Lpyki3, Zoyki3, Noyki3, 1'b0}; 
assign Juski3 = (E0yki3[3:0] | B6ski3); 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Vxyki3 
if (Dwrki3 == 1'b0) begin 
Oxyki3 <= 1'b0; 
end 
else begin 
Oxyki3 <= R1tki3; 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Hyyki3 
if (Dwrki3 == 1'b0) begin 
Cwyki3 <= 1'b0; 
end 
else begin 
Cwyki3 <= Sgski3; 
end 
end 
always @(posedge Yvrki3 or negedge Dwrki3) begin : Uyyki3 
if (Dwrki3 == 1'b0) begin 
Uzxki3 <= {32 {1'b0}}; 
end 
else 
begin 
if (Rvyki3 == 1'b1) begin 
Uzxki3 <= W1tki3; 
end 
else 
begin 
if (O8yki3 == 1'b1) begin 
Uzxki3 <= (Uzxki3 - 1); 
end 
end 
end 
end 
endmodule 
module ahb_wrapper(bus_hbusreq, bus_hgrant, bus_hlock, hsel, hclk, hresetn, pause,  
haddr_m1, hburst_m1, hbusreq_m1, hlock_m1, hprot_m1, hsize_m1, htrans_m1,  
hwdata_m1, hwrite_m1, hgrant_m1, haddr_m2, hburst_m2, hbusreq_m2, hlock_m2,  
hprot_m2, hsize_m2, htrans_m2, hwdata_m2, hwrite_m2, hgrant_m2, haddr_m3,  
hburst_m3, hbusreq_m3, hlock_m3, hprot_m3, hsize_m3, htrans_m3, hwdata_m3,  
hwrite_m3, hgrant_m3, hsel_s1, hready_resp_s1, hresp_s1, hrdata_s1, hsel_s2,  
hready_resp_s2, hresp_s2, hrdata_s2, hsplit_s2, haddr, hburst, hprot, hsize,  
htrans, hwdata, hwrite, hready, hresp, hrdata, ahbarbint, hmaster, hmaster_data, 
hmastlock); 
parameter Jsski3 = 32; 
parameter Xyrki3 = 32; 
parameter Vsski3 = 0; 
parameter Pcxki3 = 32'h01000000; 
parameter Zcxki3 = 32'h01ffffff; 
parameter Jdxki3 = 32'h02000000; 
parameter Tdxki3 = 32'h02ffffff; 
parameter Dltki3 = 128; 
parameter Rltki3 = 128; 
parameter Fmtki3 = 96; 
output [(4 - 1):0] hsel; 
output [3:0] bus_hbusreq; 
output [3:0] bus_hlock; 
output [3:0] bus_hgrant; 
input hclk; 
input hresetn; 
input pause; 
input [(Jsski3 - 1):0] haddr_m1; 
input hbusreq_m1; 
input [(3 - 1):0] hburst_m1; 
input hlock_m1; 
input [(4 - 1):0] hprot_m1; 
input [(3 - 1):0] hsize_m1; 
input [(2 - 1):0] htrans_m1; 
input [(Xyrki3 - 1):0] hwdata_m1; 
input hwrite_m1; 
output hgrant_m1; 
input [(Jsski3 - 1):0] haddr_m2; 
input hbusreq_m2; 
input [(3 - 1):0] hburst_m2; 
input hlock_m2; 
input [(4 - 1):0] hprot_m2; 
input [(3 - 1):0] hsize_m2; 
input [(2 - 1):0] htrans_m2; 
input [(Xyrki3 - 1):0] hwdata_m2; 
input hwrite_m2; 
output hgrant_m2; 
input [(Jsski3 - 1):0] haddr_m3; 
input hbusreq_m3; 
input [(3 - 1):0] hburst_m3; 
input hlock_m3; 
input [(4 - 1):0] hprot_m3; 
input [(3 - 1):0] hsize_m3; 
input [(2 - 1):0] htrans_m3; 
input [(Xyrki3 - 1):0] hwdata_m3; 
input hwrite_m3; 
output hgrant_m3; 
input hready_resp_s1; 
input [(2 - 1):0] hresp_s1; 
input [(Xyrki3 - 1):0] hrdata_s1; 
output hsel_s1; 
input hready_resp_s2; 
input [(2 - 1):0] hresp_s2; 
input [(Xyrki3 - 1):0] hrdata_s2; 
input [(16 - 1):0] hsplit_s2; 
output hsel_s2; 
output [(Jsski3 - 1):0] haddr; 
output [(3 - 1):0] hburst; 
output [(4 - 1):0] hprot; 
output [(3 - 1):0] hsize; 
output [(2 - 1):0] htrans; 
output [(Xyrki3 - 1):0] hwdata; 
output hwrite; 
output [(4 - 1):0] hmaster; 
output [(4 - 1):0] hmaster_data; 
output hmastlock; 
output ahbarbint; 
output hready; 
output [(2 - 1):0] hresp; 
output [(Xyrki3 - 1):0] hrdata; 
wire Ygski3; 
wire Hcxki3; 
wire Zdski3; 
wire [(Dltki3 - 1):0] Ogtki3; 
wire [(8 - 1):0] Ditki3; 
wire [2:0] Eezki3; 
wire [(32 - 1):0] J3ski3; 
wire [(6 - 1):0] Vjtki3; 
wire [(3 - 1):0] Kjtki3; 
wire [(Fmtki3 - 1):0] Fktki3; 
wire [(12 - 1):0] Ygtki3; 
wire [(12 - 1):0] Thtki3; 
wire [(16 - 1):0] Jhtki3; 
wire [(4 - 1):0] Zitki3; 
wire [(Rltki3 - 1):0] Oitki3; 
wire Nezki3; 
wire Iiski3; 
wire [(Xyrki3 - 1):0] Gjski3; 
wire [(2 - 1):0] Xiski3; 
wire Zwrki3; 
wire [(2 - 1):0] Ayrki3; 
wire Jxrki3; 
wire [(Xyrki3 - 1):0] Lyrki3; 
wire Vezki3; 
wire Ffzki3; 
wire Ufzki3; 
wire Ggzki3; 
wire [3:1] Mrski3; 
wire Yrski3; 
wire [(32 - 1):0] Zgzki3; 
wire [(32 - 1):0] Qhzki3; 
wire [(32 - 1):0] Hizki3; 
wire [(32 - 1):0] Yizki3; 
wire [(32 - 1):0] Pjzki3; 
wire [(32 - 1):0] Gkzki3; 
wire [(32 - 1):0] Xkzki3; 
wire [(32 - 1):0] Nlzki3; 
wire [(32 - 1):0] Dmzki3; 
wire [(32 - 1):0] Tmzki3; 
wire [(32 - 1):0] Jnzki3; 
wire [(32 - 1):0] Znzki3; 
wire [(32 - 1):0] Pozki3; 
wire [(32 - 1):0] Fpzki3; 
wire [(32 - 1):0] Vpzki3; 
assign Ogtki3[(Jsski3 - 1):0] = {Jsski3 {1'b0}}; 
assign Ditki3[(2 - 1):0] = 2'b0; 
assign Oitki3[(Xyrki3 - 1):0] = {Xyrki3 {1'b0}}; 
assign Thtki3[(3 - 1):0] = 3'b0; 
assign Ygtki3[(3 - 1):0] = 3'b0; 
assign Jhtki3[(4 - 1):0] = 4'h3; 
assign Zitki3[0] = 1'b0; 
assign Ogtki3[((Jsski3 * 2) - 1):(Jsski3 * 1)] = haddr_m1; 
assign Ditki3[3:2] = htrans_m1; 
assign Ygtki3[5:3] = hburst_m1; 
assign Thtki3[5:3] = hsize_m1; 
assign Jhtki3[7:4] = hprot_m1; 
assign Zitki3[1] = hwrite_m1; 
assign Oitki3[((Xyrki3 * 2) - 1):(Xyrki3 * 1)] = hwdata_m1; 
assign bus_hbusreq[1] = hbusreq_m1; 
assign hgrant_m1 = bus_hgrant[1]; 
assign bus_hlock[1] = hlock_m1; 
assign Ogtki3[((Jsski3 * 3) - 1):(Jsski3 * 2)] = haddr_m2; 
assign Ditki3[5:4] = htrans_m2; 
assign Ygtki3[8:6] = hburst_m2; 
assign Thtki3[8:6] = hsize_m2; 
assign Jhtki3[11:8] = hprot_m2; 
assign Zitki3[2] = hwrite_m2; 
assign Oitki3[((Xyrki3 * 3) - 1):(Xyrki3 * 2)] = hwdata_m2; 
assign bus_hbusreq[2] = hbusreq_m2; 
assign hgrant_m2 = bus_hgrant[2]; 
assign bus_hlock[2] = hlock_m2; 
assign Ogtki3[((Jsski3 * 4) - 1):(Jsski3 * 3)] = haddr_m3; 
assign Ditki3[7:6] = htrans_m3; 
assign Ygtki3[11:9] = hburst_m3; 
assign Thtki3[11:9] = hsize_m3; 
assign Jhtki3[15:12] = hprot_m3; 
assign Zitki3[3] = hwrite_m3; 
assign Oitki3[((Xyrki3 * 4) - 1):(Xyrki3 * 3)] = hwdata_m3; 
assign bus_hbusreq[3] = hbusreq_m3; 
assign hgrant_m3 = bus_hgrant[3]; 
assign bus_hlock[3] = hlock_m3; 
assign bus_hbusreq[0] = 1'b0; 
assign bus_hlock[0] = 1'b0; 
assign Kjtki3[0] = Iiski3; 
assign Vjtki3[1:0] = Xiski3; 
assign Fktki3[(Xyrki3 - 1):0] = Gjski3; 
assign Kjtki3[1] = hready_resp_s1; 
assign Vjtki3[3:2] = hresp_s1; 
assign Fktki3[((Xyrki3 * 2) - 1):(Xyrki3 * 1)] = hrdata_s1; 
assign Kjtki3[2] = hready_resp_s2; 
assign Vjtki3[5:4] = hresp_s2; 
assign Fktki3[((Xyrki3 * 3) - 1):(Xyrki3 * 2)] = hrdata_s2; 
assign Zwrki3 = hsel[(2 + 1)]; 
assign Nezki3 = hsel[0]; 
assign hsel_s1 = hsel[1]; 
assign hsel_s2 = hsel[2]; 
assign Eezki3 = hsel[2:0]; 
assign J3ski3[15:0] = {16 {1'b0}}; 
assign J3ski3[31:16] = hsplit_s2; 
assign Ufzki3 = ((0 == 1'b1) ? Hcxki3 : 1'b1); 
assign Ggzki3 = ((0 == 1'b1) ? Ygski3 : 1'b1); 
assign Vezki3 = ((1 == 1'b1) ? pause : 1'b0); 
assign Ffzki3 = ((1'b0 == 1'b1) ? Zdski3 : 1'b0); 
Dgtki3 #(Jsski3, Xyrki3) Lqzki3( .Yvrki3 (hclk),  .Dwrki3 (hresetn),  .Ogtki3 
(Ogtki3),  .Ygtki3 (Ygtki3),  .Qjski3 (hmaster),  .Jhtki3 (Jhtki3),  .Thtki3 
(Thtki3),  .Ditki3 (Ditki3),  .Oitki3 (Oitki3),  .Zitki3 (Zitki3),  .Lyrki3 
(Lyrki3),  .Jxrki3 (Jxrki3),  .Ayrki3 (Ayrki3),  .Kjtki3 (Kjtki3),  .Vjtki3 
(Vjtki3),  .Fktki3 (Fktki3),  .Keski3 (hsel[2:0]),  .U3ski3 (hmaster_data),  
.Peski3 (haddr),  .Veski3 (hburst),  .Qktki3 (hprot),  .Cfski3 (hsize),  .Swrki3 
(htrans),  .Ifski3 (hwdata),  .Pfski3 (hwrite),  .Wktki3 (hrdata),  .Lwrki3 
(hready),  .D3ski3 (hresp)); 
Vbxki3 #(Jsski3, Pcxki3, Zcxki3, Jdxki3, Tdxki3) Rqzki3( .Peski3 (haddr),  
.Hcxki3 (Ufzki3),  .Keski3 (hsel)); 
Odski3 #(Jsski3, Xyrki3, Vsski3) Yqzki3( .Yvrki3 (hclk),  .Dwrki3 (hresetn),  
.Zdski3 (Ffzki3),  .Lwrki3 (hready),  .D3ski3 (hresp),  .Keski3 (Nezki3),  
.Peski3 (haddr),  .Veski3 (hburst),  .Cfski3 (hsize),  .Swrki3 (htrans),  
.Ifski3 (hwdata),  .Pfski3 (hwrite),  .Wfski3 (bus_hlock),  .Ggski3 
(bus_hbusreq),  .J3ski3 (J3ski3),  .U3ski3 (hmaster_data),  .Sgski3 (Vezki3),  
.Ygski3 (Ggzki3),  .Nhski3 (bus_hgrant),  .Yhski3 (ahbarbint),  .Iiski3 
(Iiski3),  .Xiski3 (Xiski3),  .Gjski3 (Gjski3),  .Qjski3 (hmaster),  .Yjski3 
(hmastlock),  .Ikski3 (Zgzki3),  .Vkski3 (Qhzki3),  .Ilski3 (Hizki3),  .Vlski3 
(Yizki3),  .Imski3 (Pjzki3),  .Vmski3 (Gkzki3),  .Inski3 (Xkzki3),  .Unski3 
(Nlzki3),  .Goski3 (Dmzki3),  .Soski3 (Tmzki3),  .Epski3 (Jnzki3),  .Qpski3 
(Znzki3),  .Cqski3 (Pozki3),  .Oqski3 (Fpzki3),  .Arski3 (Vpzki3),  .Mrski3 
(Mrski3),  .Yrski3 (Yrski3)); 
Jvrki3 #(Xyrki3) Erzki3( .Yvrki3 (hclk),  .Dwrki3 (hresetn),  .Lwrki3 (hready),  
.Swrki3 (htrans),  .Zwrki3 (Zwrki3),  .Jxrki3 (Jxrki3),  .Ayrki3 (Ayrki3),  
.Lyrki3 (Lyrki3)); 
endmodule 
module F6tki3(C7tki3, G7tki3, M7tki3, U7tki3, D8tki3, B6ski3, Ewski3, I8tki3,  
Azski3, Tuski3, Q8tki3); 
parameter V9ski3 = 4; 
parameter Orzki3 = 2; 
parameter Wrzki3 = 1; 
parameter Gszki3 = 0; 
parameter Rszki3 = 1; 
input C7tki3; 
input G7tki3; 
input [(V9ski3 - 1):0] M7tki3; 
input [(V9ski3 - 1):0] D8tki3; 
input [(V9ski3 - 1):0] B6ski3; 
input [((Orzki3 * V9ski3) - 1):0] U7tki3; 
output Ewski3; 
output I8tki3; 
output Azski3; 
output [(V9ski3 - 1):0] Tuski3; 
output [(((V9ski3 > 16) ? ((V9ski3 > 64) ? ((V9ski3 > 128) ? 8 : 7) : ((V9ski3 > 
32) ? 6 : 5)) : ((V9ski3 > 4) ? ((V9ski3 > 8) ? 4 : 3) : ((V9ski3 > 2) ? 2 : 1)) 
) - 1):0] Q8tki3; 
integer Muzki3; 
integer Cvzki3; 
reg Tvzki3; 
reg Fwzki3; 
reg Rwzki3; 
reg Exzki3; 
reg Qxzki3; 
reg Byzki3; 
reg [(V9ski3 - 1):0] Myzki3; 
reg Dzzki3; 
reg Mzzki3; 
reg Wzzki3; 
reg F00li3; 
reg P00li3; 
reg W00li3; 
reg D10li3; 
reg [((Orzki3 * V9ski3) - 1):0] O10li3; 
integer G30li3; 
integer U30li3; 
integer P9ski3; 
integer Dtzki3[(V9ski3 - 1):0]; 
integer Utzki3[(V9ski3 - 1):0]; 
integer B20li3[(V9ski3 - 1):0]; 
integer R20li3[(V9ski3 - 1):0]; 
event O40li3; 
event J50li3; 
assign Tuski3 = ((Muzki3 == (-2)) ? {V9ski3 {1'bx}} : (((Cvzki3 == (-1)) && ( 
Rszki3 == 0)) ? {V9ski3 {1'b0}} : ((Rszki3 == 0) ? (1'b1 << Cvzki3) : (1'b1 <<  
Muzki3)))); 
assign Q8tki3 = ((Muzki3 == (-2)) ? {((V9ski3 > 16) ? ((V9ski3 > 64) ? ((V9ski3  
> 128) ? 8 : 7) : ((V9ski3 > 32) ? 6 : 5)) : ((V9ski3 > 4) ? ((V9ski3 > 8) ? 4 : 
3) : ((V9ski3 > 2) ? 2 : 1))) {1'bx}} : (((Muzki3 == (-1)) && (Rszki3 == 1)) ? { 
((V9ski3 > 16) ? ((V9ski3 > 64) ? ((V9ski3 > 128) ? 8 : 7) : ((V9ski3 > 32) ? 6 
: 5)) : ((V9ski3 > 4) ? ((V9ski3 > 8) ? 4 : 3) : ((V9ski3 > 2) ? 2 : 1))) {1'b1} 
} : (((Cvzki3 == (-1)) && (Rszki3 == 0)) ? {((V9ski3 > 16) ? ((V9ski3 > 64) ? (( 
V9ski3 > 128) ? 8 : 7) : ((V9ski3 > 32) ? 6 : 5)) : ((V9ski3 > 4) ? ((V9ski3 > 8 
) ? 4 : 3) : ((V9ski3 > 2) ? 2 : 1))) {1'b1}} : ((Rszki3 == 0) ?  
Cvzki3[(((V9ski3 > 16) ? ((V9ski3 > 64) ? ((V9ski3 > 128) ? 8 : 7) : ((V9ski3 > 
32) ? 6 : 5)) : ((V9ski3 > 4) ? ((V9ski3 > 8) ? 4 : 3) : ((V9ski3 > 2) ? 2 : 
1))) - 1):0] : Muzki3[(((V9ski3 > 16) ? ((V9ski3 > 64) ? ((V9ski3 > 128) ? 8 : 
7) : ((V9ski3 > 32) ? 6 : 5)) : ((V9ski3 > 4) ? ((V9ski3 > 8) ? 4 : 3) : 
((V9ski3 > 2) ? 2 : 1))) - 1):0])))); 
assign I8tki3 = ((Rszki3 == 0) ? Rwzki3 : Fwzki3); 
assign Ewski3 = ((Rszki3 == 0) ? Tvzki3 : Qxzki3); 
assign Azski3 = ((Rszki3 == 0) ? Exzki3 : Byzki3); 
always @(Muzki3 or Fwzki3 or M7tki3 or D8tki3 or B6ski3 or U7tki3 or J50li3)  
begin : C60li3 
F00li3 = (^M7tki3); 
P00li3 = (^D8tki3); 
W00li3 = (^B6ski3); 
D10li3 = (^U7tki3); 
G30li3 = (-1); 
Dzzki3 = 1'b0; 
Mzzki3 = 1'b0; 
Wzzki3 = 1'b0; 
for (P9ski3 = 0; (P9ski3 < V9ski3); P9ski3 = (P9ski3 + 1)) 
R20li3[P9ski3] = Dtzki3[P9ski3]; 
U30li3 = 0; 
O10li3 = U7tki3; 
for (P9ski3 = 0; (P9ski3 < V9ski3); P9ski3 = (P9ski3 + 1)) begin 
B20li3[P9ski3] = O10li3[(Orzki3 - 1):0]; 
O10li3 = (O10li3 >> Orzki3); 
end 
Myzki3 = (M7tki3 & (~B6ski3)); 
if ((Muzki3 < (-1)) && (D8tki3 !== {V9ski3 {1'b0}})) begin 
G30li3 = (-2); 
Wzzki3 = 1'bx; 
Mzzki3 = 1'bx; 
end 
else if ((Muzki3 >= 0) && (D8tki3[Muzki3] !== 1'b0)) begin 
if (D8tki3[Muzki3] === 1'b1) begin 
G30li3 = Muzki3; 
Wzzki3 = 1'b1; 
Mzzki3 = 1'b1; 
if (Fwzki3 === 1'b0) begin 
U30li3 = 1; 
end 
end 
else 
begin 
G30li3 = (-2); 
Wzzki3 = 1'bx; 
Mzzki3 = 1'bx; 
Dzzki3 = 1'b0; 
end 
end 
else if (Myzki3 !== {V9ski3 {1'b0}}) begin 
if ((F00li3 === 1'bx) || (D10li3 === 1'bx)) begin 
G30li3 = (-2); 
Mzzki3 = 1'bx; 
Dzzki3 = 1'bx; 
end 
else 
begin 
for (P9ski3 = 0; (P9ski3 < V9ski3); P9ski3 = (P9ski3 + 1)) begin 
if (Myzki3[P9ski3] === 1'b1) begin 
if ((G30li3 < 0) || ((B20li3[P9ski3] < B20li3[G30li3]) || ((B20li3[P9ski3] ==  
B20li3[G30li3]) && (Dtzki3[P9ski3] < Dtzki3[G30li3])))) begin 
G30li3 = P9ski3; 
Mzzki3 = 1'b1; 
end 
end 
end 
U30li3 = 1; 
end 
end 
else if (Wrzki3 == 1) begin 
G30li3 = Gszki3; 
Dzzki3 = 1'b1; 
end 
else 
begin 
G30li3 = (-1); 
end 
for (P9ski3 = 0; (P9ski3 < V9ski3); P9ski3 = (P9ski3 + 1)) begin 
if (P9ski3 == G30li3) begin 
R20li3[P9ski3] = ((1 << ((V9ski3 > 16) ? ((V9ski3 > 64) ? ((V9ski3 > 128) ? 8 :  
7) : ((V9ski3 > 32) ? 6 : 5)) : ((V9ski3 > 4) ? ((V9ski3 > 8) ? 4 : 3) : (( 
V9ski3 > 2) ? 2 : 1)))) - 1); 
end 
else if (Myzki3[P9ski3] == 1'b1) begin 
if (U30li3 == 1) begin 
if (R20li3[P9ski3] == 0) begin 
R20li3[P9ski3] = ((1 << ((V9ski3 > 16) ? ((V9ski3 > 64) ? ((V9ski3 > 128) ? 8 :  
7) : ((V9ski3 > 32) ? 6 : 5)) : ((V9ski3 > 4) ? ((V9ski3 > 8) ? 4 : 3) : (( 
V9ski3 > 2) ? 2 : 1)))) - 1); 
end 
else begin 
R20li3[P9ski3] = (Dtzki3[P9ski3] - 1); 
end 
end 
end 
else 
begin 
R20li3[P9ski3] = ((1 << ((V9ski3 > 16) ? ((V9ski3 > 64) ? ((V9ski3 > 128) ? 8 :  
7) : ((V9ski3 > 32) ? 6 : 5)) : ((V9ski3 > 4) ? ((V9ski3 > 8) ? 4 : 3) : (( 
V9ski3 > 2) ? 2 : 1)))) - 1); 
end 
end 
Cvzki3 = G30li3; 
Tvzki3 = Dzzki3; 
Rwzki3 = Mzzki3; 
Exzki3 = Wzzki3; 
for (P9ski3 = 0; (P9ski3 < V9ski3); P9ski3 = (P9ski3 + 1)) 
Utzki3[P9ski3] = R20li3[P9ski3]; 
end 
always @(posedge C7tki3 or negedge G7tki3) begin : R60li3 
if (G7tki3 === 1'b0) begin 
Muzki3 <= (-1); 
Qxzki3 <= 1'b0; 
Fwzki3 <= 1'b0; 
Byzki3 <= 1'b0; 
for (P9ski3 = 0; (P9ski3 < V9ski3); P9ski3 = (P9ski3 + 1)) 
Dtzki3[P9ski3] <= ((1 << ((V9ski3 > 16) ? ((V9ski3 > 64) ? ((V9ski3 > 128) ? 8 : 
7) : ((V9ski3 > 32) ? 6 : 5)) : ((V9ski3 > 4) ? ((V9ski3 > 8) ? 4 : 3) : (( 
V9ski3 > 2) ? 2 : 1)))) - 1); 
-> O40li3; 
end 
else if (G7tki3 === 1'b1) begin 
Muzki3 <= Cvzki3; 
Qxzki3 <= Tvzki3; 
Fwzki3 <= Rwzki3; 
Byzki3 <= Exzki3; 
for (P9ski3 = 0; (P9ski3 < V9ski3); P9ski3 = (P9ski3 + 1)) begin 
if (Dtzki3[P9ski3] !== Utzki3[P9ski3]) begin 
Dtzki3[P9ski3] <= Utzki3[P9ski3]; 
-> O40li3; 
end 
end 
end 
else 
begin 
Muzki3 <= (-2); 
Qxzki3 <= 1'bx; 
Fwzki3 <= 1'bx; 
Byzki3 <= 1'bx; 
for (P9ski3 = 0; (P9ski3 < V9ski3); P9ski3 = (P9ski3 + 1)) begin 
if (Dtzki3[P9ski3] !== (-1)) begin 
Dtzki3[P9ski3] <= (-1); 
-> O40li3; 
end 
end 
end 
end 
always @(O40li3) begin : F70li3 
#(1) ; 
-> J50li3; 
end 
initial begin : Z70li3 
integer P80li3; 
P80li3 = 0; 
if ((V9ski3 < 2) || (V9ski3 > 32)) begin 
P80li3 = 1; 
$display( 
"ERROR: %m :\n  Invalid value (%d) for parameter n (legal range: 2 to 32)",  
V9ski3); 
end 
if ((Orzki3 < 1) || (Orzki3 > 5)) begin 
P80li3 = 1; 
$display( 
"ERROR: %m :\n  Invalid value (%d) for parameter p_width (legal range: 1 to 5)", 
Orzki3); 
end 
if ((Wrzki3 < 0) || (Wrzki3 > 1)) begin 
P80li3 = 1; 
$display( 
"ERROR: %m :\n  Invalid value (%d) for parameter park_mode (legal range: 0 to 1)", 
Wrzki3); 
end 
if ((Gszki3 < 0) || (Gszki3 > (V9ski3 - 1))) begin 
P80li3 = 1; 
$display( 
"ERROR: %m :\n  Invalid value (%d) for parameter park_index (legal range: 0 to n-1)", 
Gszki3); 
end 
if ((Rszki3 < 0) || (Rszki3 > 1)) begin 
P80li3 = 1; 
$display( 
"ERROR: %m :\n  Invalid value (%d) for parameter output_mode (legal range: 0 to 1)", 
Rszki3); 
end 
if (P80li3 == 1) begin 
$display("%m :\n  Simulation aborted due to invalid parameter value(s)"); 
$finish; 
end 
end 
always @(C7tki3) begin : U90li3 
if (((C7tki3 !== 1'b0) && (C7tki3 !== 1'b1)) && ($time > 0)) begin 
$display( 
"WARNING: %m :\n  at time = %t, detected unknown value, %b, on clk input.",  
$time, C7tki3); 
end 
end 
endmodule 
module Tntki3(Kotki3, Motki3, Qotki3); 
parameter Ma0li3 = 8; 
parameter Ua0li3 = 2; 
parameter Eb0li3 = 2; 
input [(Ma0li3 - 1):0] Kotki3; 
input [(Ua0li3 - 1):0] Motki3; 
output [(Eb0li3 - 1):0] Qotki3; 
assign Qotki3[(Eb0li3 - 1):0] = (((^(Motki3 ^ Motki3)) !== 1'b0) ? {Eb0li3 {1'bx 
}} : Ob0li3(Kotki3, Motki3)); 
function [(Eb0li3 - 1):0] Ob0li3; 
input [(Ma0li3 - 1):0] Wb0li3; 
input [(Ua0li3 - 1):0] Yb0li3; 
reg [(Ma0li3 - 1):0] Wb0li3; 
reg [(Ua0li3 - 1):0] Yb0li3; 
integer P9ski3; 
integer R9ski3; 
reg [(Eb0li3 - 1):0] Cc0li3; 
begin 
for (P9ski3 = 0; (P9ski3 < Eb0li3); P9ski3 = (P9ski3 + 1)) begin 
R9ski3 = ((Yb0li3 * Eb0li3) + P9ski3); 
if (R9ski3 > (Ma0li3 - 1)) begin 
Cc0li3[P9ski3] = 1'b0; 
end 
else begin 
Cc0li3[P9ski3] = Wb0li3[R9ski3]; 
end 
end 
Ob0li3 = Cc0li3; 
end 
endfunction 
initial begin : Z70li3 
integer P80li3; 
P80li3 = 0; 
if (Ma0li3 < 1) begin 
P80li3 = 1; 
$display( 
"ERROR: %m :\n  Invalid value (%d) for parameter A_width (lower bound: 1)",  
Ma0li3); 
end 
if (Ua0li3 < 1) begin 
P80li3 = 1; 
$display( 
"ERROR: %m :\n  Invalid value (%d) for parameter SEL_width (lower bound: 1)",  
Ua0li3); 
end 
if (Eb0li3 < 1) begin 
P80li3 = 1; 
$display( 
"ERROR: %m :\n  Invalid value (%d) for parameter MUX_width (lower bound: 1)",  
Eb0li3); 
end 
if (P80li3 == 1) begin 
$display("%m :\n  Simulation aborted due to invalid parameter value(s)"); 
$finish; 
end 
end 
endmodule 
