module Fd0dwq2(Ud0dwq2,Zd0dwq2,He0dwq2,Oe0dwq2,Ve0dwq2,Ff0dwq2,Wf0dwq2,
Hg0dwq2);input Ud0dwq2;
input Zd0dwq2;
input He0dwq2;
input[(2-1):0]Oe0dwq2;
input Ve0dwq2;
output Ff0dwq2;
output[(2-1):0]Wf0dwq2;
`define L3lkc `AHB_DATA_WIDTH
output[(`L3lkc-1):0]Hg0dwq2;
reg Ff0dwq2;
reg[(2-1):0]Wf0dwq2;
reg Tg0dwq2;
reg Hh0dwq2;
wire Sh0dwq2;assign Sh0dwq2=(((Oe0dwq2==2'b11)||(Oe0dwq2==2'b10))&&((Ve0dwq2==1'b1)&&(He0dwq2==1'b1)));assign Hg0dwq2={`L3lkc {1'b0}};
always @(Tg0dwq2 or Sh0dwq2)begin : Fi0dwq2 case(Tg0dwq2)1'b0: begin if(Sh0dwq2==1'b1)begin Hh0dwq2=1'b1;end else begin Hh0dwq2=1'b0;
end end default: begin Hh0dwq2=1'b0;end endcase end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Vi0dwq2 if(Zd0dwq2==1'b0)begin 
Tg0dwq2 <=1'b0;end else begin Tg0dwq2 <=Hh0dwq2;end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Oj0dwq2 if(Zd0dwq2==1'b0)begin 
Ff0dwq2 <=1'b1;Wf0dwq2 <=2'b0;end else begin case(Tg0dwq2)1'b0: begin if(Sh0dwq2==1'b1)begin Ff0dwq2 <=1'b0;Wf0dwq2 <=2'b1;
end else begin Ff0dwq2 <=1'b1;Wf0dwq2 <=2'b0;end end default: begin Ff0dwq2 <=1'b1;Wf0dwq2 <=2'b1;end endcase end end endmodule 
module Yj0dwq2(Ud0dwq2,Zd0dwq2,Kk0dwq2,Qk0dwq2,Bl0dwq2,Ol0dwq2,Zl0dwq2,Mm0dwq2,He0dwq2,Rm0dwq2,Ym0dwq2);input Ud0dwq2;
input Zd0dwq2;input[(2-1):0]Kk0dwq2;input[(32-1):0]Qk0dwq2;input[(4-1):0]Bl0dwq2;input Mm0dwq2;input[1:0]Ol0dwq2;
input[((4*2)-1):0]Zl0dwq2;input He0dwq2;output[(16-1):0]Rm0dwq2;output[1:0]Ym0dwq2;reg[(16-1):0]Rm0dwq2;reg[1:0]Ym0dwq2;
reg[(32-1):0]Dn0dwq2;reg[(16-1):0]Qn0dwq2;reg[(2-1):0]Bo0dwq2;reg[3:0]No0dwq2;reg[3:0]Yo0dwq2;integer Op0dwq2;
integer Qp0dwq2;integer Sp0dwq2;integer Up0dwq2;integer Wp0dwq2;integer Yp0dwq2;always @(Qk0dwq2)begin : Aq0dwq2 for(Sp0dwq2=0;(Sp0dwq2 <=(16-1));Sp0dwq2=(Sp0dwq2+1))begin 
for(Up0dwq2=0;(Up0dwq2 < 2);Up0dwq2=(Up0dwq2+1))begin Dn0dwq2[((Sp0dwq2*2)+Up0dwq2)]=Qk0dwq2[((16*Up0dwq2)+Sp0dwq2)];
end end end always @(Dn0dwq2)begin : Rq0dwq2 Rm0dwq2={16 {1'b0}};for(Wp0dwq2=0;(Wp0dwq2 <=(16-1));Wp0dwq2=(Wp0dwq2+1))begin 
Bo0dwq2=(Dn0dwq2 >>(2*Wp0dwq2));Rm0dwq2[Wp0dwq2]=(|Bo0dwq2);end end always @(Kk0dwq2 or Qn0dwq2 or Rm0dwq2 or Bl0dwq2 or Zl0dwq2 or Mm0dwq2 or  
He0dwq2 or Ol0dwq2)begin : Dr0dwq2 Ym0dwq2=16'b0;case(Bl0dwq2)4'b0: Yp0dwq2=0;4'b1: Yp0dwq2=4;4'h2: Yp0dwq2=8;4'h3: 
Yp0dwq2=12;4'h4: Yp0dwq2=16;4'h5: Yp0dwq2=20;4'h6: Yp0dwq2=24;4'h7: Yp0dwq2=28;4'h8: Yp0dwq2=32;4'h9: Yp0dwq2=36;
4'ha: Yp0dwq2=40;4'hb: Yp0dwq2=44;4'hc: Yp0dwq2=48;4'hd: Yp0dwq2=52;4'he: Yp0dwq2=56;4'hf: Yp0dwq2=60;default: Yp0dwq2=0;
endcase Yo0dwq2=(Zl0dwq2 >> Yp0dwq2);for(Op0dwq2=0;(Op0dwq2 < 2);Op0dwq2=(Op0dwq2+1))begin No0dwq2=(Zl0dwq2 >>(4*Op0dwq2));
Ym0dwq2[Op0dwq2]=(((((Ol0dwq2[Op0dwq2]==1'b1)||(((Kk0dwq2==2'b11)&&(Bl0dwq2==Op0dwq2))&&(He0dwq2==1'b0)))||((Qn0dwq2[Op0dwq2]==1'b1)&&(
Rm0dwq2[Op0dwq2]==1'b0)))||((((Mm0dwq2==1'b0)&&(Kk0dwq2==2'b10))&&(No0dwq2 > Yo0dwq2))&&(He0dwq2==1'b0)))||((((Mm0dwq2==1'b1)&&(Kk0dwq2  
==2'b10))&&(Bl0dwq2 !=Op0dwq2))&&(He0dwq2==1'b0)));end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Nr0dwq2 if(Zd0dwq2==1'b0)begin 
Qn0dwq2 <={16 {1'b0}};end else begin for(Qp0dwq2=0;(Qp0dwq2 < 16);Qp0dwq2=(Qp0dwq2+1))begin if(((Kk0dwq2==2'b11)&&(He0dwq2==1'b0))&&(Bl0dwq2==Qp0dwq2))begin 
Qn0dwq2[Qp0dwq2]<=1'b1;end else begin if(Rm0dwq2[Qp0dwq2]==1'b1)begin Qn0dwq2[Qp0dwq2]<=1'b0;end end end end end endmodule 
module Ds0dwq2(Ud0dwq2,Zd0dwq2,He0dwq2,Kk0dwq2,Os0dwq2,Ts0dwq2,Zs0dwq2,Gt0dwq2,Oe0dwq2,Mt0dwq2,Tt0dwq2,Au0dwq2,Ku0dwq2,Qk0dwq2,Bl0dwq2,Wu0dwq2,
Cv0dwq2,Nv0dwq2,Xv0dwq2,Mw0dwq2,Vw0dwq2,Fx0dwq2,Nx0dwq2,Xx0dwq2,Jy0dwq2);input Ud0dwq2;input Zd0dwq2;input He0dwq2;input[(2-1):0]Kk0dwq2;
input Os0dwq2;input[(32-1):0]Ts0dwq2;input[(3-1):0]Zs0dwq2;input[(3-1):0]Gt0dwq2;input[(2-1):0]Oe0dwq2;input[(`L3lkc-1):0]Mt0dwq2;
input Tt0dwq2;input[1:0]Au0dwq2;input[1:0]Ku0dwq2;input[(32-1):0]Qk0dwq2;input[(4-1):0]Bl0dwq2;input Wu0dwq2;output[1:0]Cv0dwq2;
output Nv0dwq2;output Xv0dwq2;output[(2-1):0]Mw0dwq2;output[(`L3lkc-1):0]Vw0dwq2;output[(4-1):0]Fx0dwq2;output Nx0dwq2;
output[1:1]Xx0dwq2;output Jy0dwq2;wire Uy0dwq2;wire[((4*2)-1):0]Zl0dwq2;wire[(16-1):0]Rm0dwq2;wire[9:0]Gz0dwq2;
wire[(4-1):0]Pz0dwq2;wire[1:0]Ol0dwq2;wire[1:0]Ym0dwq2;wire[1:0]Xz0dwq2;wire[1:0]H01dwq2;wire[1:0]N01dwq2;wire[1:0]W01dwq2;
wire F11dwq2;wire M11dwq2;wire W11dwq2;wire G21dwq2;wire M21dwq2;wire X21dwq2;wire F31dwq2;wire N31dwq2;reg[255:0]U31dwq2;
wire F41dwq2;wire T41dwq2;wire[1:0]F51dwq2;wire[(480-1):0]S51dwq2;wire E61dwq2;wire[(32-1):0]J61dwq2;wire Mm0dwq2;
assign Xx0dwq2[1]=((0==1)? Xz0dwq2[1]: {1 {1'b0}});assign Jy0dwq2=((0==1)? Uy0dwq2 : 1'b0);assign X21dwq2=((1==0)? 1'b0 : T41dwq2);
assign Nv0dwq2=((1==0)? 1'b0 : F41dwq2);S61dwq2 F71dwq2(.Ud0dwq2(Ud0dwq2),.Zd0dwq2(Zd0dwq2),.Os0dwq2(Os0dwq2),.He0dwq2(He0dwq2),.Fx0dwq2(Fx0dwq2),.X21dwq2(X21dwq2),.Ts0dwq2 
(Ts0dwq2),.Oe0dwq2(Oe0dwq2),.Gt0dwq2(Gt0dwq2),.Mt0dwq2(U31dwq2),.Tt0dwq2(Tt0dwq2),.Xv0dwq2(Xv0dwq2),.Mw0dwq2(Mw0dwq2),.Vw0dwq2 
(Vw0dwq2),.M21dwq2(M21dwq2),.Gz0dwq2(Gz0dwq2),.G21dwq2(G21dwq2),.Pz0dwq2(Pz0dwq2),.Zl0dwq2(Zl0dwq2),.Ol0dwq2(Ol0dwq2),.E61dwq2 
(E61dwq2),.S51dwq2(S51dwq2),.J61dwq2(J61dwq2));C81dwq2 N81dwq2(.Ud0dwq2(Ud0dwq2),.Zd0dwq2(Zd0dwq2),.Gz0dwq2(Gz0dwq2),
.G21dwq2(G21dwq2),.M21dwq2(M21dwq2),.He0dwq2(He0dwq2),.F31dwq2(F31dwq2),.Nv0dwq2(F41dwq2),.X21dwq2(T41dwq2));Yj0dwq2 T81dwq2(.Ud0dwq2(Ud0dwq2),.Zd0dwq2(Zd0dwq2),.Kk0dwq2(Kk0dwq2),
.Qk0dwq2(Qk0dwq2),.Bl0dwq2(Bl0dwq2),.Ol0dwq2(Ol0dwq2),.Zl0dwq2(Zl0dwq2),.Mm0dwq2(Mm0dwq2),.He0dwq2(He0dwq2),.Rm0dwq2(Rm0dwq2),
.Ym0dwq2(Ym0dwq2));A91dwq2 N91dwq2(.Ud0dwq2(Ud0dwq2),.Zd0dwq2(Zd0dwq2),.Au0dwq2(Au0dwq2),.Pz0dwq2(Pz0dwq2),.Wu0dwq2(Wu0dwq2),.Zs0dwq2(Zs0dwq2),.He0dwq2 
(He0dwq2),.Kk0dwq2(Kk0dwq2),.Rm0dwq2(Rm0dwq2),.Oe0dwq2(Oe0dwq2),.N01dwq2(N01dwq2),.M11dwq2(M11dwq2),.Ym0dwq2(Ym0dwq2),.X21dwq2 
(X21dwq2),.Mm0dwq2(Mm0dwq2),.Ku0dwq2(Ku0dwq2),.F51dwq2(F51dwq2),.Cv0dwq2(Cv0dwq2),.Nx0dwq2(Nx0dwq2),.Fx0dwq2(Fx0dwq2),.F31dwq2 
(F31dwq2));V91dwq2 #(2,4,1,0,0)Ja1dwq2(.Sa1dwq2(Ud0dwq2),.Wa1dwq2(Zd0dwq2),.Cb1dwq2(F51dwq2),.Kb1dwq2(Zl0dwq2),.Tb1dwq2({(1+1){1'b0}}),.Ym0dwq2 
(Ym0dwq2),.F11dwq2(F11dwq2),.H01dwq2(H01dwq2));V91dwq2 #(2,4,1,0,0)Sc1dwq2(.Sa1dwq2(Ud0dwq2),.Wa1dwq2(Zd0dwq2),.Cb1dwq2(F51dwq2),.Kb1dwq2(Zl0dwq2),.Tb1dwq2({(1+1){1'b0}}),.Ym0dwq2 
(Xz0dwq2),.F11dwq2(W11dwq2),.H01dwq2(W01dwq2));Bd1dwq2 Pd1dwq2(.E61dwq2(E61dwq2),.N01dwq2(N01dwq2),.M11dwq2(M11dwq2),
.H01dwq2(H01dwq2),.F11dwq2(F11dwq2),.W01dwq2(W01dwq2),.W11dwq2(W11dwq2));always @(Mt0dwq2)begin : N71dwq2 U31dwq2=256'b0;
U31dwq2[(`L3lkc-1):0]=Mt0dwq2;end endmodule module C81dwq2(Ud0dwq2,Zd0dwq2,He0dwq2,Gz0dwq2,G21dwq2,M21dwq2,F31dwq2,Nv0dwq2,X21dwq2);
parameter Yd1dwq2=2'b0;parameter Ae1dwq2=2'b1;parameter Ce1dwq2=2'b11;input Ud0dwq2;input Zd0dwq2;input He0dwq2;input[9:0]Gz0dwq2;
input G21dwq2;input M21dwq2;input F31dwq2;output Nv0dwq2;output X21dwq2;reg[9:0]Ee1dwq2;wire[9:0]Oe1dwq2;reg F41dwq2;reg Ue1dwq2;
reg Hf1dwq2;wire Xf1dwq2;reg[1:0]Jg1dwq2;wire[1:0]Tg0dwq2;reg[1:0]Hh0dwq2;assign Tg0dwq2=((1==1'b1)? Jg1dwq2 : Yd1dwq2);
assign Oe1dwq2=((1==1'b1)? Ee1dwq2 : 10'b0);assign Nv0dwq2=((1==1'b1)? F41dwq2 : 1'b0);assign Xf1dwq2=((1==1'b1)? Hf1dwq2 : 1'b0);
assign X21dwq2=(Ue1dwq2 | Xf1dwq2);always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Bh1dwq2 if(Zd0dwq2==1'b0)begin Jg1dwq2 <=Yd1dwq2;
end else begin Jg1dwq2 <=Hh0dwq2;end end always @(Tg0dwq2 or G21dwq2 or F31dwq2 or Oe1dwq2)begin : Fi0dwq2 case(Tg0dwq2)Yd1dwq2: begin 
if((G21dwq2==1'b1)&&(F31dwq2==1'b1))begin Hh0dwq2=Ae1dwq2;end else begin Hh0dwq2=Yd1dwq2;end end Ae1dwq2: begin if(G21dwq2==1'b1)begin 
if(F31dwq2==1'b1)begin Hh0dwq2=Ae1dwq2;end else begin if(Oe1dwq2==10'b1)begin Hh0dwq2=Ce1dwq2;end else begin Hh0dwq2=Ae1dwq2;
end end end else begin Hh0dwq2=Yd1dwq2;end end Ce1dwq2: begin if(G21dwq2==1'b1)begin if(F31dwq2==1'b1)begin Hh0dwq2=Ae1dwq2;
end else begin Hh0dwq2=Yd1dwq2;end end else begin Hh0dwq2=Yd1dwq2;end end default: Hh0dwq2=Yd1dwq2;endcase end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Th1dwq2 
if(Zd0dwq2==1'b0)begin Ee1dwq2 <=10'b0;end else begin if(Tg0dwq2==Ce1dwq2)begin Ee1dwq2 <=Gz0dwq2;end else begin if(F31dwq2==1'b1)begin 
Ee1dwq2 <=Gz0dwq2;end else begin Ee1dwq2 <=(Ee1dwq2-10'b1);end end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Ei1dwq2 
if(Zd0dwq2==1'b0)begin F41dwq2 <=1'b0;end else begin if(G21dwq2==1'b0)begin F41dwq2 <=1'b0;end else begin if((X21dwq2==1'b1)&&(He0dwq2==1'b1))begin 
F41dwq2 <=1'b1;end else begin if(M21dwq2==1'b1)begin F41dwq2 <=1'b0;end end end end end always @(Tg0dwq2 or G21dwq2)begin : Ti1dwq2 
if(Tg0dwq2==Ce1dwq2)begin Ue1dwq2=G21dwq2;end else begin Ue1dwq2=1'b0;end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Lj1dwq2 
if(Zd0dwq2==1'b0)begin Hf1dwq2 <=1'b0;end else begin if(G21dwq2==1'b1)begin if(He0dwq2==1'b0)begin if(Ue1dwq2==1'b1)begin 
Hf1dwq2 <=1'b1;end end else begin Hf1dwq2 <=1'b0;end end else begin Hf1dwq2 <=1'b0;end end end endmodule module Ck1dwq2(Ud0dwq2,Zd0dwq2,Nk1dwq2,Xk1dwq2,Fx0dwq2,Il1dwq2,Sl1dwq2,
Cm1dwq2,Nm1dwq2,Ym1dwq2,Hg0dwq2,Ff0dwq2,Wf0dwq2,Jn1dwq2,Un1dwq2,Eo1dwq2,Os0dwq2,Bl0dwq2,Ts0dwq2,Zs0dwq2,Po1dwq2,Gt0dwq2,Oe0dwq2,Mt0dwq2,Tt0dwq2,
Vo1dwq2,He0dwq2,Kk0dwq2);input Ud0dwq2;input Zd0dwq2;input[(((1+1)*32)-1):0]Nk1dwq2;input[(6-1):0]Xk1dwq2;input[(4-1):0]Fx0dwq2;
input[(8-1):0]Il1dwq2;input[(6-1):0]Sl1dwq2;input[(4-1):0]Cm1dwq2;input[((2*`L3lkc)-1):0]Nm1dwq2;input[(2-1):0]Ym1dwq2;
input[(`L3lkc-1):0]Hg0dwq2;input[((3*`L3lkc)-1):0]Eo1dwq2;input Ff0dwq2;input[(2-1):0]Wf0dwq2;input[(3-1):0]Jn1dwq2;
input[(6-1):0]Un1dwq2;input[2:0]Os0dwq2;output[(32-1):0]Ts0dwq2;output[(3-1):0]Zs0dwq2;output[(4-1):0]Po1dwq2;
output[(3-1):0]Gt0dwq2;output[(2-1):0]Oe0dwq2;output[(`L3lkc-1):0]Mt0dwq2;output Tt0dwq2;output[(4-1):0]Bl0dwq2;
output[(`L3lkc-1):0]Vo1dwq2;output He0dwq2;output[(2-1):0]Kk0dwq2;reg[(4-1):0]Bl0dwq2;reg[(`L3lkc-1):0]Vo1dwq2;
reg He0dwq2;reg[(2-1):0]Kk0dwq2;reg[2:0]Cp1dwq2;integer Qp0dwq2;Mp1dwq2 #(((1+1)*32),4,32)Zp1dwq2(.Dq1dwq2(Nk1dwq2),.Fq1dwq2 
(Fx0dwq2),.Jq1dwq2(Ts0dwq2));Mp1dwq2 #(4,4,2)Nq1dwq2(.Dq1dwq2(Cm1dwq2),.Fq1dwq2(Fx0dwq2),.Jq1dwq2(Oe0dwq2));Mp1dwq2 #(6,4,3)Rq1dwq2(.Dq1dwq2(Xk1dwq2),.Fq1dwq2(Fx0dwq2),.Jq1dwq2 
(Zs0dwq2));Mp1dwq2 #(6,4,3)Vq1dwq2(.Dq1dwq2(Sl1dwq2),.Fq1dwq2(Fx0dwq2),.Jq1dwq2(Gt0dwq2));Mp1dwq2 #(8,4,4)Zq1dwq2(.Dq1dwq2(Il1dwq2),.Fq1dwq2(Fx0dwq2),.Jq1dwq2 
(Po1dwq2));Mp1dwq2 #(2,4,1)Dr1dwq2(.Dq1dwq2(Ym1dwq2),.Fq1dwq2(Fx0dwq2),.Jq1dwq2(Tt0dwq2));Mp1dwq2 #((2*`L3lkc),4,`L3lkc)Ir1dwq2(.Dq1dwq2(Nm1dwq2),.Fq1dwq2(Bl0dwq2),
.Jq1dwq2(Mt0dwq2));always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Nr1dwq2 if(Zd0dwq2==1'b0)begin Bl0dwq2 <={4 {1'b0}};
end else begin if(He0dwq2==1'b1)begin Bl0dwq2 <=Fx0dwq2;end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Fs1dwq2 
if(Zd0dwq2==1'b0)begin Cp1dwq2 <={(2+1){1'b0}};end else begin if(He0dwq2==1'b1)begin Cp1dwq2 <=Os0dwq2;end end end always @(Cp1dwq2 or Eo1dwq2 or Jn1dwq2 or Un1dwq2 or Wf0dwq2 or Hg0dwq2 or  
Ff0dwq2)begin : Us1dwq2 He0dwq2=Ff0dwq2;Kk0dwq2=Wf0dwq2;Vo1dwq2=Hg0dwq2;for(Qp0dwq2=0;(Qp0dwq2 <=2);Qp0dwq2=(Qp0dwq2+1))begin 
if(Cp1dwq2[Qp0dwq2]==1'b1)begin He0dwq2=Jn1dwq2[Qp0dwq2];Kk0dwq2=(Un1dwq2 >>(Qp0dwq2*2));Vo1dwq2=(Eo1dwq2 >>(Qp0dwq2*`L3lkc));
end end end endmodule module S61dwq2(Ud0dwq2,Zd0dwq2,Os0dwq2,He0dwq2,Fx0dwq2,X21dwq2,Ts0dwq2,Oe0dwq2,Gt0dwq2,Mt0dwq2,Tt0dwq2,Xv0dwq2,Mw0dwq2,Vw0dwq2,M21dwq2,Gz0dwq2,
G21dwq2,Pz0dwq2,Zl0dwq2,Ol0dwq2,E61dwq2,S51dwq2,J61dwq2);parameter Hb2dwq2=2'b0;parameter Pb2dwq2=2'b1;parameter Xb2dwq2=2'b10;
parameter Gc2dwq2=2'b11;input Ud0dwq2;input Zd0dwq2;input Os0dwq2;input He0dwq2;input[(32-1):0]Ts0dwq2;input[(2-1):0]Oe0dwq2;
input[(3-1):0]Gt0dwq2;input[255:0]Mt0dwq2;input Tt0dwq2;input[(4-1):0]Fx0dwq2;input X21dwq2;output Xv0dwq2;output[(2-1):0]Mw0dwq2;
output[(`L3lkc-1):0]Vw0dwq2;output[9:0]Gz0dwq2;output G21dwq2;output[(4-1):0]Pz0dwq2;output M21dwq2;output[((4*2)-1):0]Zl0dwq2;
output[1:0]Ol0dwq2;output E61dwq2;output[(480-1):0]S51dwq2;output[(32-1):0]J61dwq2;reg M21dwq2;wire Sh0dwq2;wire Qt1dwq2;
wire Au1dwq2;wire Ku1dwq2;wire Su1dwq2;wire Av1dwq2;wire Iv1dwq2;wire Qv1dwq2;wire Yv1dwq2;wire Gw1dwq2;wire Ow1dwq2;wire Ww1dwq2;
wire Ex1dwq2;wire Nx1dwq2;wire Wx1dwq2;wire Fy1dwq2;wire Oy1dwq2;wire Xy1dwq2;wire Gz1dwq2;wire Tz1dwq2;wire D02dwq2;wire P02dwq2;
wire[255:0]T02dwq2;wire[15:0]H12dwq2;wire[63:0]W12dwq2;wire[3:0]N22dwq2;wire[3:0]X22dwq2;wire[3:0]H32dwq2;wire[3:0]R32dwq2;
wire[3:0]B42dwq2;wire[3:0]L42dwq2;wire[3:0]V42dwq2;wire[3:0]F52dwq2;wire[3:0]P52dwq2;wire[3:0]Z52dwq2;wire[3:0]K62dwq2;
wire[3:0]V62dwq2;wire[3:0]G72dwq2;wire[3:0]R72dwq2;wire[3:0]C82dwq2;wire[9:0]N82dwq2;wire[9:0]X82dwq2;wire[(4-1):0]M92dwq2;
wire Z92dwq2;wire Ja2dwq2;wire Va2dwq2;reg[3:0]Pc2dwq2;reg[3:0]Uc2dwq2;reg[3:0]Zc2dwq2;reg[3:0]Ed2dwq2;reg[3:0]Jd2dwq2;
reg[3:0]Od2dwq2;reg[3:0]Td2dwq2;reg[3:0]Yd2dwq2;reg[3:0]De2dwq2;reg[3:0]Ie2dwq2;reg[3:0]Oe2dwq2;reg[3:0]Ue2dwq2;
reg[3:0]Af2dwq2;reg[3:0]Gf2dwq2;reg[3:0]Mf2dwq2;wire[3:0]Sf2dwq2;wire[3:0]Wf2dwq2;wire[3:0]Ag2dwq2;wire[3:0]Eg2dwq2;
wire[3:0]Ig2dwq2;wire[3:0]Mg2dwq2;wire[3:0]Qg2dwq2;wire[3:0]Ug2dwq2;wire[3:0]Yg2dwq2;wire[3:0]Ch2dwq2;wire[3:0]Hh2dwq2;
wire[3:0]Mh2dwq2;wire[3:0]Rh2dwq2;wire[3:0]Wh2dwq2;wire[3:0]Bi2dwq2;reg[9:0]Gi2dwq2;reg Qi2dwq2;reg[3:0]Xi2dwq2;
reg Gj2dwq2;reg Xj2dwq2;reg[(2-1):0]Nk2dwq2;reg Yk2dwq2;reg Jl2dwq2;reg[(4-1):0]Wl2dwq2;reg[(32-1):0]Im2dwq2;reg[(2-1):0]Sm2dwq2;
reg[(3-1):0]Dn2dwq2;wire[(32-1):0]Nn2dwq2;wire[(2-1):0]Vn2dwq2;wire[(3-1):0]Eo2dwq2;wire Mo2dwq2;wire Vo2dwq2;
wire[(4-1):0]Gp2dwq2;reg[1:0]Qp2dwq2;wire[1:0]Yp2dwq2;reg[1:0]Eq2dwq2;reg[31:0]Oq2dwq2;reg[31:0]Zq2dwq2;reg[31:0]Hr2dwq2;
reg Tr2dwq2;wire Bs2dwq2;reg Fs2dwq2;wire[(32-1):0]Rs2dwq2;wire[(32-1):0]Gt2dwq2;wire[(32-1):0]Vt2dwq2;wire[(32-1):0]Ku2dwq2;
wire[(32-1):0]Zu2dwq2;wire[(32-1):0]Ov2dwq2;wire[(32-1):0]Dw2dwq2;wire[(32-1):0]Sw2dwq2;wire[(32-1):0]Hx2dwq2;
wire[(32-1):0]Wx2dwq2;wire[(32-1):0]My2dwq2;wire[(32-1):0]Cz2dwq2;wire[(32-1):0]Sz2dwq2;wire[(32-1):0]I03dwq2;
wire[(32-1):0]Y03dwq2;reg O13dwq2;wire U13dwq2;wire F23dwq2;reg[31:0]O23dwq2;reg[31:0]E33dwq2;reg[31:0]U33dwq2;reg[31:0]K43dwq2;
reg[31:0]A53dwq2;reg[31:0]Q53dwq2;reg[31:0]G63dwq2;reg[31:0]W63dwq2;reg[31:0]M73dwq2;reg[31:0]C83dwq2;reg[31:0]T83dwq2;
reg[31:0]K93dwq2;reg[31:0]Ba3dwq2;reg[31:0]Sa3dwq2;reg[31:0]Jb3dwq2;wire[(32-1):0]Ac3dwq2;wire[(32-1):0]Oc3dwq2;
reg[(32-1):0]Yc3dwq2;reg[31:0]Hd3dwq2;wire Td3dwq2;reg[(32-1):0]Fe3dwq2;reg[(32-1):0]Re3dwq2;reg[(32-1):0]Df3dwq2;
reg[(32-1):0]Pf3dwq2;reg[(32-1):0]Bg3dwq2;reg[(32-1):0]Ng3dwq2;reg[(32-1):0]Zg3dwq2;reg[(32-1):0]Lh3dwq2;reg[(32-1):0]Xh3dwq2;
reg[(32-1):0]Ji3dwq2;reg[(32-1):0]Wi3dwq2;reg[(32-1):0]Jj3dwq2;reg[(32-1):0]Wj3dwq2;reg[(32-1):0]Jk3dwq2;reg[(32-1):0]Wk3dwq2;
wire[(32-1):0]Jl3dwq2;wire[(32-1):0]Wl3dwq2;wire[(32-1):0]Jm3dwq2;wire[(32-1):0]Wm3dwq2;wire[(32-1):0]Jn3dwq2;
wire[(32-1):0]Wn3dwq2;wire[(32-1):0]Jo3dwq2;wire[(32-1):0]Wo3dwq2;wire[(32-1):0]Jp3dwq2;wire[(32-1):0]Wp3dwq2;
wire[(32-1):0]Kq3dwq2;wire[(32-1):0]Yq3dwq2;wire[(32-1):0]Mr3dwq2;wire[(32-1):0]As3dwq2;wire[(32-1):0]Os3dwq2;
wire[(32-1):0]Ct3dwq2;wire[(32-1):0]Tt3dwq2;wire[(32-1):0]Ku3dwq2;wire[(32-1):0]Bv3dwq2;wire[(32-1):0]Sv3dwq2;
wire[(32-1):0]Jw3dwq2;wire[(32-1):0]Ax3dwq2;wire[(32-1):0]Rx3dwq2;wire[(32-1):0]Iy3dwq2;wire[(32-1):0]Zy3dwq2;
wire[(32-1):0]Rz3dwq2;wire[(32-1):0]J04dwq2;wire[(32-1):0]B14dwq2;wire[(32-1):0]T14dwq2;wire[(32-1):0]L24dwq2;
wire D34dwq2;wire O34dwq2;wire Z34dwq2;wire K44dwq2;wire V44dwq2;wire G54dwq2;wire R54dwq2;wire C64dwq2;wire N64dwq2;wire Y64dwq2;
wire K74dwq2;wire W74dwq2;wire I84dwq2;wire U84dwq2;wire G94dwq2;assign Sh0dwq2=((Oe0dwq2 !=2'b0)&&(Oe0dwq2 !=2'b1));assign Qt1dwq2=((Os0dwq2==1'b1)&&(He0dwq2==1'b1));
assign Au1dwq2=((Qt1dwq2==1'b1)&&(Sh0dwq2==1'b1));assign Vo2dwq2=((1==1)? Jl2dwq2 : 1'b0);assign Mo2dwq2=((1==1)? Yk2dwq2 : 1'b0);
assign Nn2dwq2=((1==1)? Im2dwq2 : {32 {1'b0}});assign Vn2dwq2=((1==1)? Sm2dwq2 : {2 {1'b0}});assign Eo2dwq2=((1==1)? Dn2dwq2 : {4 {1'b0}});
assign Gp2dwq2=((1==1)? Wl2dwq2 : {4 {1'b0}});assign Z92dwq2=((Vn2dwq2 !=2'b0)&&(Vn2dwq2 !=2'b1));assign Ja2dwq2=((Z92dwq2==1'b1)&&(Vo2dwq2==1'b1));
assign Mw0dwq2=((1==1'b1)? Nk2dwq2 : {2 {1'b0}});assign Xv0dwq2=((1==1'b1)? Gj2dwq2 : 1'b1);assign Yp2dwq2=((1==1'b1)? Qp2dwq2 : Hb2dwq2);
assign P02dwq2=(((Mo2dwq2==1'b1)&&(Ja2dwq2==1'b1))&&(He0dwq2==1'b1));assign Ku1dwq2=((Nn2dwq2[9:0]==10'b0)&&(P02dwq2==1'b1));
assign Su1dwq2=((Nn2dwq2[9:0]==10'h004)&&(P02dwq2==1'b1));assign Av1dwq2=((Nn2dwq2[9:0]==10'h008)&&(P02dwq2==1'b1));
assign Iv1dwq2=((Nn2dwq2[9:0]==10'h00c)&&(P02dwq2==1'b1));assign Qv1dwq2=((Nn2dwq2[9:0]==10'h010)&&(P02dwq2==1'b1));
assign Yv1dwq2=((Nn2dwq2[9:0]==10'h014)&&(P02dwq2==1'b1));assign Gw1dwq2=((Nn2dwq2[9:0]==10'h018)&&(P02dwq2==1'b1));
assign Ow1dwq2=((Nn2dwq2[9:0]==10'h01c)&&(P02dwq2==1'b1));assign Ww1dwq2=((Nn2dwq2[9:0]==10'h020)&&(P02dwq2==1'b1));
assign Ex1dwq2=((Nn2dwq2[9:0]==10'h024)&&(P02dwq2==1'b1));assign Nx1dwq2=((Nn2dwq2[9:0]==10'h028)&&(P02dwq2==1'b1));
assign Wx1dwq2=((Nn2dwq2[9:0]==10'h02c)&&(P02dwq2==1'b1));assign Fy1dwq2=((Nn2dwq2[9:0]==10'h030)&&(P02dwq2==1'b1));
assign Oy1dwq2=((Nn2dwq2[9:0]==10'h034)&&(P02dwq2==1'b1));assign Xy1dwq2=((Nn2dwq2[9:0]==10'h038)&&(P02dwq2==1'b1));
assign Gz1dwq2=((Nn2dwq2[9:0]==10'h03c)&&(P02dwq2==1'b1));assign Tz1dwq2=((Nn2dwq2[9:0]==10'h040)&&(P02dwq2==1'b1));
assign D02dwq2=((Nn2dwq2[9:0]==10'h048)&&(P02dwq2==1'b1));assign F23dwq2=((Nn2dwq2[9:0]==10'h04c)&&(P02dwq2==1'b1));
assign Td3dwq2=((Nn2dwq2[9:0]==10'h050)&&(P02dwq2==1'b1));assign D34dwq2=((Nn2dwq2[9:0]==10'h054)&&(P02dwq2==1'b1));
assign O34dwq2=((Nn2dwq2[9:0]==10'h058)&&(P02dwq2==1'b1));assign Z34dwq2=((Nn2dwq2[9:0]==10'h05c)&&(P02dwq2==1'b1));
assign K44dwq2=((Nn2dwq2[9:0]==10'h060)&&(P02dwq2==1'b1));assign V44dwq2=((Nn2dwq2[9:0]==10'h064)&&(P02dwq2==1'b1));
assign G54dwq2=((Nn2dwq2[9:0]==10'h068)&&(P02dwq2==1'b1));assign R54dwq2=((Nn2dwq2[9:0]==10'h06c)&&(P02dwq2==1'b1));
assign C64dwq2=((Nn2dwq2[9:0]==10'h070)&&(P02dwq2==1'b1));assign N64dwq2=((Nn2dwq2[9:0]==10'h074)&&(P02dwq2==1'b1));
assign Y64dwq2=((Nn2dwq2[9:0]==10'h078)&&(P02dwq2==1'b1));assign K74dwq2=((Nn2dwq2[9:0]==10'h07c)&&(P02dwq2==1'b1));
assign W74dwq2=((Nn2dwq2[9:0]==10'h080)&&(P02dwq2==1'b1));assign I84dwq2=((Nn2dwq2[9:0]==10'h084)&&(P02dwq2==1'b1));
assign U84dwq2=((Nn2dwq2[9:0]==10'h088)&&(P02dwq2==1'b1));assign G94dwq2=((Nn2dwq2[9:0]==10'h08c)&&(P02dwq2==1'b1));
assign N22dwq2=Oq2dwq2[3:0];assign Sf2dwq2=(((1==0)||(0==1))? 4'b1 : Pc2dwq2);assign X22dwq2=Oq2dwq2[3:0];assign Wf2dwq2=((1 < 2)? 4'b0 :(((1==0)||(0==1))? 4'h2 : Uc2dwq2));
assign H32dwq2=Oq2dwq2[3:0];assign Ag2dwq2=((1 < 3)? 4'b0 :(((1==0)||(0==1))? 4'h3 : Zc2dwq2));assign R32dwq2=Oq2dwq2[3:0];
assign Eg2dwq2=((1 < 4)? 4'b0 :(((1==0)||(0==1))? 4'h4 : Ed2dwq2));assign B42dwq2=Oq2dwq2[3:0];assign Ig2dwq2=((1 < 5)? 4'b0 :(((1==0)||(0==1))? 4'h5 : Jd2dwq2));
assign L42dwq2=Oq2dwq2[3:0];assign Mg2dwq2=((1 < 6)? 4'b0 :(((1==0)||(0==1))? 4'h6 : Od2dwq2));assign V42dwq2=Oq2dwq2[3:0];
assign Qg2dwq2=((1 < 7)? 4'b0 :(((1==0)||(0==1))? 4'h7 : Td2dwq2));assign F52dwq2=Oq2dwq2[3:0];assign Ug2dwq2=((1 < 8)? 4'b0 :(((1==0)||(0==1))? 4'h8 : Yd2dwq2));
assign P52dwq2=Oq2dwq2[3:0];assign Yg2dwq2=((1 < 9)? 4'b0 :(((1==0)||(0==1))? 4'h9 : De2dwq2));assign Z52dwq2=Oq2dwq2[3:0];
assign Ch2dwq2=((1 < 10)? 4'b0 :(((1==0)||(0==1))? 4'ha : Ie2dwq2));assign K62dwq2=Oq2dwq2[3:0];assign Hh2dwq2=((1 < 11)? 4'b0 :(((1==0)||(0==1))? 4'hb : Oe2dwq2));
assign V62dwq2=Oq2dwq2[3:0];assign Mh2dwq2=((1 < 12)? 4'b0 :(((1==0)||(0==1))? 4'hc : Ue2dwq2));assign G72dwq2=Oq2dwq2[3:0];
assign Rh2dwq2=((1 < 13)? 4'b0 :(((1==0)||(0==1))? 4'hd : Af2dwq2));assign R72dwq2=Oq2dwq2[3:0];assign Wh2dwq2=((1 < 14)? 4'b0 :(((1==0)||(0==1))? 4'he : Gf2dwq2));
assign C82dwq2=Oq2dwq2[3:0];assign Bi2dwq2=((1 < 15)? 4'b0 :(((1==0)||(0==1))? 4'hf : Mf2dwq2));assign X82dwq2=Oq2dwq2[9:0];
assign Va2dwq2=Oq2dwq2[0];assign Gz0dwq2=(((1==1'b0)||(1==1'b0))? 10'b0 : Gi2dwq2);assign G21dwq2=(((1==1'b0)||(1==1'b0))? 1'b0 : Qi2dwq2);
assign M92dwq2=Oq2dwq2[3:0];assign Pz0dwq2=(((0==1)||(1==1'b0))? 0 : Xi2dwq2);assign Bs2dwq2=(((1==1'b1)&&(1==1'b1))? Tr2dwq2 : 1'b0);
assign U13dwq2=Oq2dwq2[0];assign E61dwq2=(((0==1'b1)&&(1==1'b1))? O13dwq2 : 1'b0);assign Ac3dwq2=Oq2dwq2[(32-1):0];
assign Oc3dwq2=(((1==1)||(1==1'b0))? 32'h0000ffff : Yc3dwq2);assign J61dwq2=Oc3dwq2;assign Ct3dwq2=Oq2dwq2[(32-1):0];
assign Jl3dwq2=(((1==1)||(1==1'b0))? 32'h0000000f : Fe3dwq2);assign Tt3dwq2=Oq2dwq2[(32-1):0];assign Wl3dwq2=(((1==1)||(1==1'b0))? 32'h0000000f : Re3dwq2);
assign Ku3dwq2=Oq2dwq2[(32-1):0];assign Jm3dwq2=(((1==1)||(1==1'b0))? 32'h0000000f : Df3dwq2);assign Bv3dwq2=Oq2dwq2[(32-1):0];
assign Wm3dwq2=(((1==1)||(1==1'b0))? 32'h0000000f : Pf3dwq2);assign Sv3dwq2=Oq2dwq2[(32-1):0];assign Jn3dwq2=(((1==1)||(1==1'b0))? 32'h0000000f : Bg3dwq2);
assign Jw3dwq2=Oq2dwq2[(32-1):0];assign Wn3dwq2=(((1==1)||(1==1'b0))? 32'h0000000f : Ng3dwq2);assign Ax3dwq2=Oq2dwq2[(32-1):0];
assign Jo3dwq2=(((1==1)||(1==1'b0))? 32'h0000000f : Zg3dwq2);assign Rx3dwq2=Oq2dwq2[(32-1):0];assign Wo3dwq2=(((1==1)||(1==1'b0))? 32'h0000000f : Lh3dwq2);
assign Iy3dwq2=Oq2dwq2[(32-1):0];assign Jp3dwq2=(((1==1)||(1==1'b0))? 32'h0000000f : Xh3dwq2);assign Zy3dwq2=Oq2dwq2[(32-1):0];
assign Wp3dwq2=(((1==1)||(1==1'b0))? 32'h0000000f : Ji3dwq2);assign Rz3dwq2=Oq2dwq2[(32-1):0];assign Kq3dwq2=(((1==1)||(1==1'b0))? 32'h0000000f : Wi3dwq2);
assign J04dwq2=Oq2dwq2[(32-1):0];assign Yq3dwq2=(((1==1)||(1==1'b0))? 32'h0000000f : Jj3dwq2);assign B14dwq2=Oq2dwq2[(32-1):0];
assign Mr3dwq2=(((1==1)||(1==1'b0))? 32'h0000000f : Wj3dwq2);assign T14dwq2=Oq2dwq2[(32-1):0];assign As3dwq2=(((1==1)||(1==1'b0))? 32'h0000000f : Jk3dwq2);
assign L24dwq2=Oq2dwq2[(32-1):0];assign Os3dwq2=(((1==1)||(1==1'b0))? 32'h0000000f : Wk3dwq2);assign N82dwq2=(Xv0dwq2 ? Ts0dwq2[9:0]: Nn2dwq2[9:0]);
`define M1lkc `BIG_ENDIAN
assign T02dwq2[31:0]=((`M1lkc==1'b0)? Zq2dwq2[31:0]: {Zq2dwq2[7:0],Zq2dwq2[15:8],Zq2dwq2[23:16],Zq2dwq2[31:24]});assign T02dwq2[63:32]=T02dwq2[31:0];
assign T02dwq2[95:64]=T02dwq2[31:0];assign T02dwq2[127:96]=T02dwq2[31:0];assign T02dwq2[159:128]=T02dwq2[31:0];assign T02dwq2[191:160]=T02dwq2[31:0];
assign T02dwq2[223:192]=T02dwq2[31:0];assign T02dwq2[255:224]=T02dwq2[31:0];assign Vw0dwq2=T02dwq2[(`L3lkc-1):0];assign H12dwq2[0]=1'b0;
assign H12dwq2[1]=(Sf2dwq2[3:0]==4'b0);assign H12dwq2[2]=((1 >=2)?(Wf2dwq2[3:0]==4'b0): 1'b0);assign H12dwq2[3]=((1 >=3)?(Ag2dwq2[3:0]==4'b0): 1'b0);
assign H12dwq2[4]=((1 >=4)?(Eg2dwq2[3:0]==4'b0): 1'b0);assign H12dwq2[5]=((1 >=5)?(Ig2dwq2[3:0]==4'b0): 1'b0);assign H12dwq2[6]=((1 >=6)?(Mg2dwq2[3:0]==4'b0): 1'b0);
assign H12dwq2[7]=((1 >=7)?(Qg2dwq2[3:0]==4'b0): 1'b0);assign H12dwq2[8]=((1 >=8)?(Ug2dwq2[3:0]==4'b0): 1'b0);assign H12dwq2[9]=((1 >=9)?(Yg2dwq2[3:0]==4'b0): 1'b0);
assign H12dwq2[10]=((1 >=10)?(Ch2dwq2[3:0]==4'b0): 1'b0);assign H12dwq2[11]=((1 >=11)?(Hh2dwq2[3:0]==4'b0): 1'b0);
assign H12dwq2[12]=((1 >=12)?(Mh2dwq2[3:0]==4'b0): 1'b0);assign H12dwq2[13]=((1 >=13)?(Rh2dwq2[3:0]==4'b0): 1'b0);
assign H12dwq2[14]=((1 >=14)?(Wh2dwq2[3:0]==4'b0): 1'b0);assign H12dwq2[15]=((1==15)?(Bi2dwq2[3:0]==4'b0): 1'b0);
assign Ol0dwq2=H12dwq2[1:0];assign W12dwq2[3:0]=4'hf;assign W12dwq2[7:4]=(~Sf2dwq2[3:0]);assign W12dwq2[11:8]=(~Wf2dwq2[3:0]);
assign W12dwq2[15:12]=(~Ag2dwq2[3:0]);assign W12dwq2[19:16]=(~Eg2dwq2[3:0]);assign W12dwq2[23:20]=(~Ig2dwq2[3:0]);assign W12dwq2[27:24]=(~Mg2dwq2[3:0]);
assign W12dwq2[31:28]=(~Qg2dwq2[3:0]);assign W12dwq2[35:32]=(~Ug2dwq2[3:0]);assign W12dwq2[39:36]=(~Yg2dwq2[3:0]);assign W12dwq2[43:40]=(~Ch2dwq2[3:0]);
assign W12dwq2[47:44]=(~Hh2dwq2[3:0]);assign W12dwq2[51:48]=(~Mh2dwq2[3:0]);assign W12dwq2[55:52]=(~Rh2dwq2[3:0]);assign W12dwq2[59:56]=(~Wh2dwq2[3:0]);
assign W12dwq2[63:60]=(~Bi2dwq2[3:0]);assign Zl0dwq2=W12dwq2[((4*2)-1):0];assign Rs2dwq2=Jl3dwq2;assign Gt2dwq2=((1 >=2)? Wl3dwq2 : {32 {1'b0}});
assign Vt2dwq2=((1 >=3)? Jm3dwq2 : {32 {1'b0}});assign Ku2dwq2=((1 >=4)? Wm3dwq2 : {32 {1'b0}});assign Zu2dwq2=((1 >=5)? Jn3dwq2 : {32 {1'b0}});
assign Ov2dwq2=((1 >=6)? Wn3dwq2 : {32 {1'b0}});assign Dw2dwq2=((1 >=7)? Jo3dwq2 : {32 {1'b0}});assign Sw2dwq2=((1 >=8)? Wo3dwq2 : {32 {1'b0}});
assign Hx2dwq2=((1 >=9)? Jp3dwq2 : {32 {1'b0}});assign Wx2dwq2=((1 >=10)? Wp3dwq2 : {32 {1'b0}});assign My2dwq2=((1 >=11)? Kq3dwq2 : {32 {1'b0}});
assign Cz2dwq2=((1 >=12)? Yq3dwq2 : {32 {1'b0}});assign Sz2dwq2=((1 >=13)? Mr3dwq2 : {32 {1'b0}});assign I03dwq2=((1 >=14)? As3dwq2 : {32 {1'b0}});
assign Y03dwq2=((1 >=15)? Os3dwq2 : {32 {1'b0}});assign S51dwq2[(32-1):0]=Rs2dwq2;assign S51dwq2[((32*2)-1):32]=Gt2dwq2;
assign S51dwq2[((32*3)-1):(32*2)]=Vt2dwq2;assign S51dwq2[((32*4)-1):(32*3)]=Ku2dwq2;assign S51dwq2[((32*5)-1):(32*4)]=Zu2dwq2;
assign S51dwq2[((32*6)-1):(32*5)]=Ov2dwq2;assign S51dwq2[((32*7)-1):(32*6)]=Dw2dwq2;assign S51dwq2[((32*8)-1):(32*7)]=Sw2dwq2;
assign S51dwq2[((32*9)-1):(32*8)]=Hx2dwq2;assign S51dwq2[((32*10)-1):(32*9)]=Wx2dwq2;assign S51dwq2[((32*11)-1):(32*10)]=My2dwq2;
assign S51dwq2[((32*12)-1):(32*11)]=Cz2dwq2;assign S51dwq2[((32*13)-1):(32*12)]=Sz2dwq2;assign S51dwq2[((32*14)-1):(32*13)]=I03dwq2;
assign S51dwq2[((32*15)-1):(32*14)]=Y03dwq2;always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : S94dwq2 if(Zd0dwq2==1'b0)begin 
Jl2dwq2 <=1'b0;end else begin if(He0dwq2==1'b1)begin Jl2dwq2 <=Os0dwq2;end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Ia4dwq2 
if(Zd0dwq2==1'b0)begin Im2dwq2 <=32'b0;Sm2dwq2 <=2'b0;Yk2dwq2 <=1'b0;Dn2dwq2 <=3'b0;Wl2dwq2 <=4'b0;end else begin if(He0dwq2==1'b1)begin 
Im2dwq2 <=Ts0dwq2;Sm2dwq2 <=Oe0dwq2;Yk2dwq2 <=Tt0dwq2;Dn2dwq2 <=Gt0dwq2;Wl2dwq2 <=Fx0dwq2;end end end always @(Ts0dwq2)begin : Qa4dwq2 
Fs2dwq2=1'b0;case(Ts0dwq2[9:0])10'b0: Fs2dwq2=1'b1;10'h004: if(1 > 1)begin Fs2dwq2=1'b1;end 10'h008: if(1 > 2)begin 
Fs2dwq2=1'b1;end 10'h00c: if(1 > 3)begin Fs2dwq2=1'b1;end 10'h010: if(1 > 4)begin Fs2dwq2=1'b1;end 10'h014: if(1 > 5)begin 
Fs2dwq2=1'b1;end 10'h018: if(1 > 6)begin Fs2dwq2=1'b1;end 10'h01c: if(1 > 7)begin Fs2dwq2=1'b1;end 10'h020: if(1 > 8)begin 
Fs2dwq2=1'b1;end 10'h024: if(1 > 9)begin Fs2dwq2=1'b1;end 10'h028: if(1 > 10)begin Fs2dwq2=1'b1;end 10'h02c: if(1 > 11)begin 
Fs2dwq2=1'b1;end 10'h030: if(1 > 12)begin Fs2dwq2=1'b1;end 10'h034: if(1 > 13)begin Fs2dwq2=1'b1;end 10'h038: if(1 > 14)begin 
Fs2dwq2=1'b1;end 10'h03c: if(1==1'b1)begin Fs2dwq2=1'b1;end 10'h040: if(1==1'b1)begin Fs2dwq2=1'b1;end 10'h044: if(1==1'b1)begin 
Fs2dwq2=1'b1;end 10'h048: Fs2dwq2=1'b1;10'h04c: if(0==1'b1)begin Fs2dwq2=1'b1;end 10'h050: if(0==1'b1)begin Fs2dwq2=1'b1;
end 10'h054: if(0==1'b1)begin Fs2dwq2=1'b1;end 10'h058: if((0==1'b1)&&(1 > 1))begin Fs2dwq2=1'b1;end 10'h05c: if((0==1'b1)&&(1 > 2))begin 
Fs2dwq2=1'b1;end 10'h060: if((0==1'b1)&&(1 > 3))begin Fs2dwq2=1'b1;end 10'h064: if((0==1'b1)&&(1 > 4))begin Fs2dwq2=1'b1;
end 10'h068: if((0==1'b1)&&(1 > 5))begin Fs2dwq2=1'b1;end 10'h06c: if((0==1'b1)&&(1 > 6))begin Fs2dwq2=1'b1;end 10'h070: 
if((0==1'b1)&&(1 > 7))begin Fs2dwq2=1'b1;end 10'h074: if((0==1'b1)&&(1 > 8))begin Fs2dwq2=1'b1;end 10'h078: if((0==1'b1)&&(1 > 9))begin 
Fs2dwq2=1'b1;end 10'h07c: if((0==1'b1)&&(1 > 10))begin Fs2dwq2=1'b1;end 10'h080: if((0==1'b1)&&(1 > 11))begin Fs2dwq2=1'b1;
end 10'h084: if((0==1'b1)&&(1 > 12))begin Fs2dwq2=1'b1;end 10'h088: if((0==1'b1)&&(1 > 13))begin Fs2dwq2=1'b1;end 
10'h08c: if((0==1'b1)&&(1 > 14))begin Fs2dwq2=1'b1;end default: Fs2dwq2=1'b0;endcase end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Hb4dwq2 
if(Zd0dwq2==1'b0)begin Nk2dwq2 <=2'b0;end else begin if((Yp2dwq2==Gc2dwq2)||(Eq2dwq2==Gc2dwq2))begin Nk2dwq2 <=2'b1;
end else begin Nk2dwq2 <=2'b0;end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Xb4dwq2 if(Zd0dwq2==1'b0)begin 
Gj2dwq2 <=1'b1;end else begin Gj2dwq2 <=Xj2dwq2;end end always @(Yp2dwq2 or Eq2dwq2 or Ts0dwq2 or Nn2dwq2)begin : Rc4dwq2 if((((Yp2dwq2==Xb2dwq2)&&(Eq2dwq2==Pb2dwq2))&&(Ts0dwq2[9:0]==
Nn2dwq2[9:0]))||(Eq2dwq2==Gc2dwq2))begin Xj2dwq2=1'b0;end else begin Xj2dwq2=1'b1;end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Md4dwq2 
if(Zd0dwq2==1'b0)begin Qp2dwq2 <=Hb2dwq2;end else begin Qp2dwq2 <=Eq2dwq2;end end always @(Yp2dwq2 or Au1dwq2 or Tt0dwq2 or Fs2dwq2 or Gt0dwq2)begin : Xd4dwq2 
case(Yp2dwq2)Hb2dwq2,Xb2dwq2,Pb2dwq2: if(Au1dwq2==1'b1)begin if((Fs2dwq2==1'b1)&&(Gt0dwq2==3'b010))begin if(Tt0dwq2==1'b1)begin 
Eq2dwq2=Xb2dwq2;end else begin Eq2dwq2=Pb2dwq2;end end else begin Eq2dwq2=Gc2dwq2;end end else begin Eq2dwq2=Hb2dwq2;end 
default: Eq2dwq2=Hb2dwq2;endcase end always @(Mt0dwq2 or Nn2dwq2)begin : Me4dwq2 if(`M1lkc==0)begin if(`L3lkc==32)begin 
Oq2dwq2=Mt0dwq2[31:0];end else if(`L3lkc==64)begin case(Nn2dwq2[2:0])3'h4: Oq2dwq2=Mt0dwq2[63:32];default: Oq2dwq2=Mt0dwq2[31:0];
endcase end else if(`L3lkc==128)begin case(Nn2dwq2[3:0])4'h4: Oq2dwq2=Mt0dwq2[63:32];4'h8: Oq2dwq2=Mt0dwq2[95:64];4'hc: 
Oq2dwq2=Mt0dwq2[127:96];default: Oq2dwq2=Mt0dwq2[31:0];endcase end else begin case(Nn2dwq2[4:0])5'h04: Oq2dwq2=Mt0dwq2[63:32];
5'h08: Oq2dwq2=Mt0dwq2[95:64];5'h0c: Oq2dwq2=Mt0dwq2[127:96];5'h10: Oq2dwq2=Mt0dwq2[159:128];5'h14: Oq2dwq2=Mt0dwq2[191:160];
5'h18: Oq2dwq2=Mt0dwq2[223:192];5'h1c: Oq2dwq2=Mt0dwq2[255:224];default: Oq2dwq2=Mt0dwq2[31:0];endcase end end else if(`L3lkc==32)begin 
Oq2dwq2[7:0]=Mt0dwq2[31:24];Oq2dwq2[15:8]=Mt0dwq2[23:16];Oq2dwq2[23:16]=Mt0dwq2[15:8];Oq2dwq2[31:24]=Mt0dwq2[7:0];end else if(`L3lkc==64)begin 
case(Nn2dwq2[2:0])3'h4: begin Oq2dwq2[7:0]=Mt0dwq2[31:24];Oq2dwq2[15:8]=Mt0dwq2[23:16];Oq2dwq2[23:16]=Mt0dwq2[15:8];Oq2dwq2[31:24]=Mt0dwq2[7:0];
end default: begin Oq2dwq2[7:0]=Mt0dwq2[63:56];Oq2dwq2[15:8]=Mt0dwq2[55:48];Oq2dwq2[23:16]=Mt0dwq2[47:40];Oq2dwq2[31:24]=Mt0dwq2[39:32];
end endcase end else if(`L3lkc==128)begin case(Nn2dwq2[3:0])4'h4: begin Oq2dwq2[7:0]=Mt0dwq2[95:88];Oq2dwq2[15:8]=Mt0dwq2[87:80];
Oq2dwq2[23:16]=Mt0dwq2[79:72];Oq2dwq2[31:24]=Mt0dwq2[71:64];end 4'h8: begin Oq2dwq2[7:0]=Mt0dwq2[63:56];Oq2dwq2[15:8]=Mt0dwq2[55:48];
Oq2dwq2[23:16]=Mt0dwq2[47:40];Oq2dwq2[31:24]=Mt0dwq2[39:32];end 4'hc: begin Oq2dwq2[7:0]=Mt0dwq2[31:24];Oq2dwq2[15:8]=Mt0dwq2[23:16];
Oq2dwq2[23:16]=Mt0dwq2[15:8];Oq2dwq2[31:24]=Mt0dwq2[7:0];end default: begin Oq2dwq2[7:0]=Mt0dwq2[127:120];Oq2dwq2[15:8]=Mt0dwq2[119:112];
Oq2dwq2[23:16]=Mt0dwq2[111:104];Oq2dwq2[31:24]=Mt0dwq2[103:96];end endcase end else begin case(Nn2dwq2[4:0])5'h04: begin Oq2dwq2[7:0]=Mt0dwq2[223:216];
Oq2dwq2[15:8]=Mt0dwq2[215:208];Oq2dwq2[23:16]=Mt0dwq2[207:200];Oq2dwq2[31:24]=Mt0dwq2[199:192];end 5'h08: begin Oq2dwq2[7:0]=Mt0dwq2[191:184];
Oq2dwq2[15:8]=Mt0dwq2[183:176];Oq2dwq2[23:16]=Mt0dwq2[175:168];Oq2dwq2[31:24]=Mt0dwq2[167:160];end 5'h0c: begin Oq2dwq2[7:0]=Mt0dwq2[159:152];
Oq2dwq2[15:8]=Mt0dwq2[151:144];Oq2dwq2[23:16]=Mt0dwq2[143:136];Oq2dwq2[31:24]=Mt0dwq2[135:128];end 5'h10: begin Oq2dwq2[7:0]=Mt0dwq2[127:120];
Oq2dwq2[15:8]=Mt0dwq2[119:112];Oq2dwq2[23:16]=Mt0dwq2[111:104];Oq2dwq2[31:24]=Mt0dwq2[103:96];end 5'h14: begin Oq2dwq2[7:0]=Mt0dwq2[95:88];
Oq2dwq2[15:8]=Mt0dwq2[87:80];Oq2dwq2[23:16]=Mt0dwq2[79:72];Oq2dwq2[31:24]=Mt0dwq2[71:64];end 5'h18: begin Oq2dwq2[7:0]=Mt0dwq2[63:56];
Oq2dwq2[15:8]=Mt0dwq2[55:48];Oq2dwq2[23:16]=Mt0dwq2[47:40];Oq2dwq2[31:24]=Mt0dwq2[39:32];end 5'h1c: begin Oq2dwq2[7:0]=Mt0dwq2[31:24];
Oq2dwq2[15:8]=Mt0dwq2[23:16];Oq2dwq2[23:16]=Mt0dwq2[15:8];Oq2dwq2[31:24]=Mt0dwq2[7:0];end default: begin Oq2dwq2[7:0]=Mt0dwq2[255:248];
Oq2dwq2[15:8]=Mt0dwq2[247:240];Oq2dwq2[23:16]=Mt0dwq2[239:232];Oq2dwq2[31:24]=Mt0dwq2[231:224];end endcase end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Cf4dwq2 
if(Zd0dwq2==1'b0)begin Pc2dwq2 <=4'b1;end else begin if(Ku1dwq2==1'b1)begin if((Gp2dwq2==4'b1)&&(N22dwq2==0))begin 
Pc2dwq2 <=Pc2dwq2;end else begin Pc2dwq2 <=N22dwq2;end end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Mf4dwq2 
if(Zd0dwq2==1'b0)begin Uc2dwq2 <=4'h2;end else begin if(Su1dwq2==1'b1)begin if((Gp2dwq2==4'h2)&&(X22dwq2==0))begin 
Uc2dwq2 <=Uc2dwq2;end else begin Uc2dwq2 <=X22dwq2;end end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Wf4dwq2 
if(Zd0dwq2==1'b0)begin Zc2dwq2 <=4'h3;end else begin if(Av1dwq2==1'b1)begin if((Gp2dwq2==4'h3)&&(H32dwq2==0))begin 
Zc2dwq2 <=Zc2dwq2;end else begin Zc2dwq2 <=H32dwq2;end end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Gg4dwq2 
if(Zd0dwq2==1'b0)begin Ed2dwq2 <=4'h4;end else begin if(Iv1dwq2==1'b1)begin if((Gp2dwq2==4'h4)&&(R32dwq2==0))begin 
Ed2dwq2 <=Ed2dwq2;end else begin Ed2dwq2 <=R32dwq2;end end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Qg4dwq2 
if(Zd0dwq2==1'b0)begin Jd2dwq2 <=4'h5;end else begin if(Qv1dwq2==1'b1)begin if((Gp2dwq2==4'h5)&&(B42dwq2==0))begin 
Jd2dwq2 <=Jd2dwq2;end else begin Jd2dwq2 <=B42dwq2;end end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Ah4dwq2 
if(Zd0dwq2==1'b0)begin Od2dwq2 <=4'h6;end else begin if(Yv1dwq2==1'b1)begin if((Gp2dwq2==4'h6)&&(L42dwq2==0))begin 
Od2dwq2 <=Od2dwq2;end else begin Od2dwq2 <=L42dwq2;end end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Kh4dwq2 
if(Zd0dwq2==1'b0)begin Td2dwq2 <=4'h7;end else begin if(Gw1dwq2==1'b1)begin if((Gp2dwq2==4'h7)&&(V42dwq2==0))begin 
Td2dwq2 <=Td2dwq2;end else begin Td2dwq2 <=V42dwq2;end end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Uh4dwq2 
if(Zd0dwq2==1'b0)begin Yd2dwq2 <=4'h8;end else begin if(Ow1dwq2==1'b1)begin if((Gp2dwq2==4'h8)&&(F52dwq2==0))begin 
Yd2dwq2 <=Yd2dwq2;end else begin Yd2dwq2 <=F52dwq2;end end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Ei4dwq2 
if(Zd0dwq2==1'b0)begin De2dwq2 <=4'h9;end else begin if(Ww1dwq2==1'b1)begin if((Gp2dwq2==4'h9)&&(P52dwq2==0))begin 
De2dwq2 <=De2dwq2;end else begin De2dwq2 <=P52dwq2;end end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Oi4dwq2 
if(Zd0dwq2==1'b0)begin Ie2dwq2 <=4'ha;end else begin if(Ex1dwq2==1'b1)begin if((Gp2dwq2==4'ha)&&(Z52dwq2==0))begin 
Ie2dwq2 <=Ie2dwq2;end else begin Ie2dwq2 <=Z52dwq2;end end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Zi4dwq2 
if(Zd0dwq2==1'b0)begin Oe2dwq2 <=4'hb;end else begin if(Nx1dwq2==1'b1)begin if((Gp2dwq2==4'hb)&&(K62dwq2==0))begin 
Oe2dwq2 <=Oe2dwq2;end else begin Oe2dwq2 <=K62dwq2;end end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Kj4dwq2 
if(Zd0dwq2==1'b0)begin Ue2dwq2 <=4'hc;end else begin if(Wx1dwq2==1'b1)begin if((Gp2dwq2==4'hc)&&(V62dwq2==0))begin 
Ue2dwq2 <=Ue2dwq2;end else begin Ue2dwq2 <=V62dwq2;end end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Vj4dwq2 
if(Zd0dwq2==1'b0)begin Af2dwq2 <=4'hd;end else begin if(Fy1dwq2==1'b1)begin if((Gp2dwq2==4'hd)&&(G72dwq2==0))begin 
Af2dwq2 <=Af2dwq2;end else begin Af2dwq2 <=G72dwq2;end end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Gk4dwq2 
if(Zd0dwq2==1'b0)begin Gf2dwq2 <=4'he;end else begin if(Oy1dwq2==1'b1)begin if((Gp2dwq2==4'he)&&(R72dwq2==0))begin 
Gf2dwq2 <=Gf2dwq2;end else begin Gf2dwq2 <=R72dwq2;end end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Rk4dwq2 
if(Zd0dwq2==1'b0)begin Mf2dwq2 <=4'hf;end else begin if(Xy1dwq2==1'b1)begin if((Gp2dwq2==4'hf)&&(C82dwq2==0))begin 
Mf2dwq2 <=Mf2dwq2;end else begin Mf2dwq2 <=C82dwq2;end end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Cl4dwq2 
if(Zd0dwq2==1'b0)begin Gi2dwq2 <=10'b0;end else begin if(Gz1dwq2==1'b1)begin Gi2dwq2 <=X82dwq2;end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Rl4dwq2 
if(Zd0dwq2==1'b0)begin Qi2dwq2 <=1'b0;end else begin if(Tz1dwq2==1'b1)begin Qi2dwq2 <=Va2dwq2;end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Dm4dwq2 
if(Zd0dwq2==1'b0)begin Xi2dwq2 <=0;end else begin if(D02dwq2==1'b1)begin if(M92dwq2 > 1)begin Xi2dwq2 <={4 {1'b0}};end 
else begin Xi2dwq2 <=M92dwq2;end end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Qm4dwq2 if(Zd0dwq2==1'b0)begin 
Tr2dwq2 <=1'b0;end else begin if(X21dwq2==1'b1)begin Tr2dwq2 <=1'b1;end else begin if(M21dwq2==1'b1)begin Tr2dwq2 <=1'b0;
end end end end always @(Ts0dwq2 or Au1dwq2 or Tt0dwq2)begin : Dn4dwq2 if(((Au1dwq2==1'b1)&&(Tt0dwq2==1'b0))&&(Ts0dwq2[9:0]==10'h044))begin 
M21dwq2=1'b1;end else begin M21dwq2=1'b0;end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Tn4dwq2 if(Zd0dwq2==1'b0)begin 
O13dwq2 <=1'b0;end else begin if(F23dwq2==1'b1)begin O13dwq2 <=U13dwq2;end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Eo4dwq2 
if(Zd0dwq2==1'b0)begin Yc3dwq2 <=32'h0000ffff;end else begin if(Td3dwq2==1'b1)begin Yc3dwq2 <=Ac3dwq2;end end end always @(Oc3dwq2)begin 
Hd3dwq2=32'b0;Hd3dwq2[(32-1):0]=Oc3dwq2;end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : So4dwq2 if(Zd0dwq2==1'b0)begin 
Fe3dwq2 <=32'h0000000f;end else begin if(D34dwq2==1'b1)begin Fe3dwq2 <=Ct3dwq2;end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Jp4dwq2 
if(Zd0dwq2==1'b0)begin Re3dwq2 <=32'h0000000f;end else begin if(O34dwq2==1'b1)begin Re3dwq2 <=Tt3dwq2;end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Aq4dwq2 
if(Zd0dwq2==1'b0)begin Df3dwq2 <=32'h0000000f;end else begin if(Z34dwq2==1'b1)begin Df3dwq2 <=Ku3dwq2;end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Rq4dwq2 
if(Zd0dwq2==1'b0)begin Pf3dwq2 <=32'h0000000f;end else begin if(K44dwq2==1'b1)begin Pf3dwq2 <=Bv3dwq2;end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Ir4dwq2 
if(Zd0dwq2==1'b0)begin Bg3dwq2 <=32'h0000000f;end else begin if(V44dwq2==1'b1)begin Bg3dwq2 <=Sv3dwq2;end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Zr4dwq2 
if(Zd0dwq2==1'b0)begin Ng3dwq2 <=32'h0000000f;end else begin if(G54dwq2==1'b1)begin Ng3dwq2 <=Jw3dwq2;end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Qs4dwq2 
if(Zd0dwq2==1'b0)begin Zg3dwq2 <=32'h0000000f;end else begin if(R54dwq2==1'b1)begin Zg3dwq2 <=Ax3dwq2;end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Ht4dwq2 
if(Zd0dwq2==1'b0)begin Lh3dwq2 <=32'h0000000f;end else begin if(C64dwq2==1'b1)begin Lh3dwq2 <=Rx3dwq2;end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Yt4dwq2 
if(Zd0dwq2==1'b0)begin Xh3dwq2 <=32'h0000000f;end else begin if(N64dwq2==1'b1)begin Xh3dwq2 <=Iy3dwq2;end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Pu4dwq2 
if(Zd0dwq2==1'b0)begin Ji3dwq2 <=32'h0000000f;end else begin if(Y64dwq2==1'b1)begin Ji3dwq2 <=Zy3dwq2;end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Hv4dwq2 
if(Zd0dwq2==1'b0)begin Wi3dwq2 <=32'h0000000f;end else begin if(K74dwq2==1'b1)begin Wi3dwq2 <=Rz3dwq2;end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Zv4dwq2 
if(Zd0dwq2==1'b0)begin Jj3dwq2 <=32'h0000000f;end else begin if(W74dwq2==1'b1)begin Jj3dwq2 <=J04dwq2;end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Rw4dwq2 
if(Zd0dwq2==1'b0)begin Wj3dwq2 <=32'h0000000f;end else begin if(I84dwq2==1'b1)begin Wj3dwq2 <=B14dwq2;end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Jx4dwq2 
if(Zd0dwq2==1'b0)begin Jk3dwq2 <=32'h0000000f;end else begin if(U84dwq2==1'b1)begin Jk3dwq2 <=T14dwq2;end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : By4dwq2 
if(Zd0dwq2==1'b0)begin Wk3dwq2 <=32'h0000000f;end else begin if(G94dwq2==1'b1)begin Wk3dwq2 <=L24dwq2;end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Ty4dwq2 
if(Zd0dwq2==1'b0)begin Hr2dwq2 <=32'b0;end else begin if((Yp2dwq2==Gc2dwq2)||(Eq2dwq2==Gc2dwq2))begin Hr2dwq2 <=32'b0;
end else begin if((((Au1dwq2==1'b1)&&(Tt0dwq2==1'b0))&&(Xj2dwq2==1'b1))||(((Ja2dwq2==1'b1)&&(Mo2dwq2==1'b0))&&(Xv0dwq2==1'b0)))begin 
case(N82dwq2)10'b0: Hr2dwq2 <={28'b0,Sf2dwq2};10'h004: Hr2dwq2 <={28'b0,Wf2dwq2};10'h008: Hr2dwq2 <={28'b0,Ag2dwq2};10'h00c: 
Hr2dwq2 <={28'b0,Eg2dwq2};10'h010: Hr2dwq2 <={28'b0,Ig2dwq2};10'h014: Hr2dwq2 <={28'b0,Mg2dwq2};10'h018: Hr2dwq2 <={28'b0,Qg2dwq2};
10'h01c: Hr2dwq2 <={28'b0,Ug2dwq2};10'h020: Hr2dwq2 <={28'b0,Yg2dwq2};10'h024: Hr2dwq2 <={28'b0,Ch2dwq2};10'h028: Hr2dwq2 <={28'b0,Hh2dwq2};
10'h02c: Hr2dwq2 <={28'b0,Mh2dwq2};10'h030: Hr2dwq2 <={28'b0,Rh2dwq2};10'h034: Hr2dwq2 <={28'b0,Wh2dwq2};10'h038: Hr2dwq2 <={28'b0,Bi2dwq2};
10'h03c: Hr2dwq2 <={22'b0,Gz0dwq2};10'h040: Hr2dwq2 <={31'b0,G21dwq2};10'h044: Hr2dwq2 <={31'b0,Bs2dwq2};10'h048: Hr2dwq2 <={24'b0,Pz0dwq2};
10'h04c: Hr2dwq2 <={31'b0,E61dwq2};10'h050: Hr2dwq2 <=Hd3dwq2;10'h054: Hr2dwq2 <=O23dwq2;10'h058: Hr2dwq2 <=E33dwq2;10'h05c: 
Hr2dwq2 <=U33dwq2;10'h060: Hr2dwq2 <=K43dwq2;10'h064: Hr2dwq2 <=A53dwq2;10'h068: Hr2dwq2 <=Q53dwq2;10'h06c: Hr2dwq2 <=G63dwq2;
10'h070: Hr2dwq2 <=W63dwq2;10'h074: Hr2dwq2 <=M73dwq2;10'h078: Hr2dwq2 <=C83dwq2;10'h07c: Hr2dwq2 <=T83dwq2;10'h080: Hr2dwq2 <=K93dwq2;
10'h084: Hr2dwq2 <=Ba3dwq2;10'h088: Hr2dwq2 <=Sa3dwq2;10'h08c: Hr2dwq2 <=Jb3dwq2;endcase end end end end always @(Hr2dwq2)begin : Kz4dwq2 
Zq2dwq2=32'b0;if(1==1)begin if(0==1'b1)begin if(32 > 10)begin Zq2dwq2[(32-1):0]=Hr2dwq2[(32-1):0];end else begin 
Zq2dwq2[9:0]=Hr2dwq2[9:0];end end else begin Zq2dwq2[9:0]=Hr2dwq2[9:0];end end end always @(Rs2dwq2)begin : Xz4dwq2 O23dwq2=32'b0;
O23dwq2[(32-1):0]=Rs2dwq2;end always @(Gt2dwq2)begin : S05dwq2 E33dwq2=32'b0;E33dwq2[(32-1):0]=Gt2dwq2;end always @(Vt2dwq2)begin : N15dwq2 
U33dwq2=32'b0;U33dwq2[(32-1):0]=Vt2dwq2;end always @(Ku2dwq2)begin : I25dwq2 K43dwq2=32'b0;K43dwq2[(32-1):0]=Ku2dwq2;
end always @(Zu2dwq2)begin : D35dwq2 A53dwq2=32'b0;A53dwq2[(32-1):0]=Zu2dwq2;end always @(Ov2dwq2)begin : Y35dwq2 Q53dwq2=32'b0;
Q53dwq2[(32-1):0]=Ov2dwq2;end always @(Dw2dwq2)begin : T45dwq2 G63dwq2=32'b0;G63dwq2[(32-1):0]=Dw2dwq2;end always @(Sw2dwq2)begin : O55dwq2 
W63dwq2=32'b0;W63dwq2[(32-1):0]=Sw2dwq2;end always @(Hx2dwq2)begin : J65dwq2 M73dwq2=32'b0;M73dwq2[(32-1):0]=Hx2dwq2;
end always @(Wx2dwq2)begin : E75dwq2 C83dwq2=32'b0;C83dwq2[(32-1):0]=Wx2dwq2;end always @(My2dwq2)begin : A85dwq2 T83dwq2=32'b0;
T83dwq2[(32-1):0]=My2dwq2;end always @(Cz2dwq2)begin : W85dwq2 K93dwq2=32'b0;K93dwq2[(32-1):0]=Cz2dwq2;end always @(Sz2dwq2)begin : S95dwq2 
Ba3dwq2=32'b0;Ba3dwq2[(32-1):0]=Sz2dwq2;end always @(I03dwq2)begin : Oa5dwq2 Sa3dwq2=32'b0;Sa3dwq2[(32-1):0]=I03dwq2;
end always @(Y03dwq2)begin : Kb5dwq2 Jb3dwq2=32'b0;Jb3dwq2[(32-1):0]=Y03dwq2;end endmodule module Bd1dwq2(E61dwq2,H01dwq2,W01dwq2,F11dwq2,W11dwq2,N01dwq2,M11dwq2);
input E61dwq2;input[1:0]H01dwq2;input[1:0]W01dwq2;input F11dwq2;input W11dwq2;output[1:0]N01dwq2;output M11dwq2;reg[1:0]N01dwq2;
reg M11dwq2;always @(E61dwq2 or W11dwq2 or W01dwq2 or H01dwq2)begin N01dwq2=H01dwq2;if(0==1)begin if((E61dwq2==1'b1)&&(W11dwq2==1'b0))begin 
N01dwq2=W01dwq2;end end end always @(E61dwq2 or W11dwq2 or F11dwq2)begin M11dwq2=F11dwq2;if(0==1)begin if(E61dwq2==1'b1)begin 
M11dwq2=(F11dwq2 && W11dwq2);end end end endmodule module Gc5dwq2(Ts0dwq2,Sc5dwq2,Os0dwq2);input[(32-1):0]Ts0dwq2;input Sc5dwq2;
`define N5lkc `R1_N_SA_0
output[(4-1):0]Os0dwq2;wire[15:0]Ad5dwq2;wire[15:0]Kd5dwq2;wire[2:0]Xd5dwq2;reg Ve0dwq2;integer Op0dwq2;assign Ad5dwq2[0]=((1==1)?((Ts0dwq2 >=`N5lkc)&&(Ts0dwq2 <=
`define R7lkc `R1_N_EA_0
`define Q5lkc `R1_N_SA_1
`define T6lkc `R1_N_EA_1
`R7lkc)): 1'b0);assign Ad5dwq2[1]=((((((((((Ts0dwq2 >=`Q5lkc)&&(Ts0dwq2 <=`T6lkc))||(((Ts0dwq2 >=32'h03000000)&&(Ts0dwq2 <=32'h0300ffff))&&(
0 >=3'b1)))||(((Ts0dwq2 >=32'h04000000)&&(Ts0dwq2 <=32'h0400ffff))&&(0  >=3'b010)))||(((Ts0dwq2 >=32'h05000000)&&(Ts0dwq2 <=32'h0500ffff))&&(0  
>=3'b011)))||(((Ts0dwq2 >=32'h06000000)&&(Ts0dwq2 <=32'h0600ffff))&&(0  >=3'h4)))||(((Ts0dwq2 >=32'h07000000)&&(Ts0dwq2 <=32'h0700ffff))&&(0 >=
3'b101)))||(((Ts0dwq2 >=32'h08000000)&&(Ts0dwq2 <=32'h0800ffff))&&(0 >=3'b110)))||(((Ts0dwq2 >=32'h09000000)&&(Ts0dwq2 <=32'h0900ffff))&&(0==
`define K8lkc `R1_N_SA_2
`define E2lkc `R1_N_EA_2
`define O2lkc `R2_N_SA_2
`define W2lkc `R2_N_EA_2
3'b111)))&&(1 !=2'b10));assign Ad5dwq2[2]=((((Ts0dwq2 >=`K8lkc)&&(Ts0dwq2 <=`E2lkc))||(((Ts0dwq2 >=`O2lkc)&&(Ts0dwq2 <=`W2lkc))&&(0==1'b1)))&& 
(1 !=2'b10));assign Ad5dwq2[3]=((((Ts0dwq2 >=32'h0c000000)&&(Ts0dwq2 <=32'h0c00ffff))||(((Ts0dwq2 >=32'h0d000000)&&(Ts0dwq2 <=32'h0d00ffff))&&(0==1'b1)))&& 
(1 !=2'b10));assign Ad5dwq2[4]=((((Ts0dwq2 >=32'h0e000000)&&(Ts0dwq2 <=32'h0e00ffff))||(((Ts0dwq2 >=32'h0f000000)&&(Ts0dwq2 <=32'h0f00ffff))&&(0==1'b1)))&& 
(1 !=2'b10));assign Ad5dwq2[5]=((((Ts0dwq2 >=32'h10000000)&&(Ts0dwq2 <=32'h1000ffff))||(((Ts0dwq2 >=32'h11000000)&&(Ts0dwq2 <=32'h1100ffff))&&(0==1'b1)))&& 
(1 !=2'b10));assign Ad5dwq2[6]=((((Ts0dwq2 >=32'h12000000)&&(Ts0dwq2 <=32'h1200ffff))||(((Ts0dwq2 >=32'h13000000)&&(Ts0dwq2 <=32'h1300ffff))&&(0==1'b1)))&& 
(1 !=2'b10));assign Ad5dwq2[7]=((((Ts0dwq2 >=32'h14000000)&&(Ts0dwq2 <=32'h1400ffff))||(((Ts0dwq2 >=32'h15000000)&&(Ts0dwq2 <=32'h1500ffff))&&(0==1'b1)))&& 
(1 !=2'b10));assign Ad5dwq2[8]=((((Ts0dwq2 >=32'h16000000)&&(Ts0dwq2 <=32'h1600ffff))||(((Ts0dwq2 >=32'h17000000)&&(Ts0dwq2 <=32'h1700ffff))&&(0==1'b1)))&& 
(1 !=2'b10));assign Ad5dwq2[9]=((((Ts0dwq2 >=32'h18000000)&&(Ts0dwq2 <=32'h1800ffff))||(((Ts0dwq2 >=32'h19000000)&&(Ts0dwq2 <=32'h1900ffff))&&(0==1'b1)))&& 
(1 !=2'b10));assign Ad5dwq2[10]=((((Ts0dwq2 >=32'h1a000000)&&(Ts0dwq2 <=32'h1a00ffff))||(((Ts0dwq2 >=32'h1b000000)&&(Ts0dwq2 <=32'h1b00ffff))&&(0==1'b1)))&& 
(1 !=2'b10));assign Ad5dwq2[11]=((((Ts0dwq2 >=32'h1c000000)&&(Ts0dwq2 <=32'h1c00ffff))||(((Ts0dwq2 >=32'h1d000000)&&(Ts0dwq2 <=32'h1d00ffff))&&(0==1'b1)))&& 
(1 !=2'b10));assign Ad5dwq2[12]=((((Ts0dwq2 >=32'h1e000000)&&(Ts0dwq2 <=32'h1e00ffff))||(((Ts0dwq2 >=32'h1f000000)&&(Ts0dwq2 <=32'h1f00ffff))&&(0==1'b1)))&& 
(1 !=2'b10));assign Ad5dwq2[13]=((((Ts0dwq2 >=32'h20000000)&&(Ts0dwq2 <=32'h2000ffff))||(((Ts0dwq2 >=32'h21000000)&&(Ts0dwq2 <=32'h2100ffff))&&(0==1'b1)))&& 
(1 !=2'b10));assign Ad5dwq2[14]=((((Ts0dwq2 >=32'h22000000)&&(Ts0dwq2 <=32'h2200ffff))||(((Ts0dwq2 >=32'h23000000)&&(Ts0dwq2 <=32'h2300ffff))&&(0==1'b1)))&& 
(1 !=2'b10));assign Ad5dwq2[15]=((((Ts0dwq2 >=32'h24000000)&&(Ts0dwq2 <=32'h2400ffff))||(((Ts0dwq2 >=32'h25000000)&&(Ts0dwq2 <=32'h2500ffff))&&(0==1'b1)))&& 
(1 !=2'b10));assign Kd5dwq2[0]=((1==1)?((Ts0dwq2 >=32'h26000000)&&(Ts0dwq2 <=32'h260003ff)): 1'b0);assign Kd5dwq2[1]=((((((((((Ts0dwq2 >=32'h27000000)&&(Ts0dwq2 <=
32'h2700ffff))||(((Ts0dwq2 >=32'h28000000)&&(Ts0dwq2 <=32'h2800ffff))&&(0 >=3'b1)))||(((Ts0dwq2 >=32'h29000000)&&(Ts0dwq2 <=32'h2900ffff))&&(0  
>=3'b010)))||(((Ts0dwq2 >=32'h2a000000)&&(Ts0dwq2 <=32'h2a00ffff))&&(0  >=3'b011)))||(((Ts0dwq2 >=32'h2b000000)&&(Ts0dwq2 <=32'h2b00ffff))&&(0  
>=3'h4)))||(((Ts0dwq2 >=32'h2c000000)&&(Ts0dwq2 <=32'h2c00ffff))&&(0 >=3'b101)))||(((Ts0dwq2 >=32'h2d000000)&&(Ts0dwq2 <=32'h2d00ffff))&&(0 >=
3'b110)))||(((Ts0dwq2 >=32'h2e000000)&&(Ts0dwq2 <=32'h2e00ffff))&&(0==3'b111)))&&(1 !=2'b1));assign Kd5dwq2[2]=((((Ts0dwq2 >=32'h2f000000)&&(Ts0dwq2 <=32'h2f00ffff))
||(((Ts0dwq2 >=32'h30000000)&&(Ts0dwq2 <=32'h3000ffff))&&(0==1'b1)))&&(1 !=2'b1));assign Kd5dwq2[3]=((((Ts0dwq2 >=32'h31000000)&&(Ts0dwq2 <=32'h3100ffff))
||(((Ts0dwq2 >=32'h32000000)&&(Ts0dwq2 <=32'h3200ffff))&&(0==1'b1)))&&(1 !=2'b1));assign Kd5dwq2[4]=((((Ts0dwq2 >=32'h33000000)&&(Ts0dwq2 <=32'h3300ffff))
||(((Ts0dwq2 >=32'h34000000)&&(Ts0dwq2 <=32'h3400ffff))&&(0==1'b1)))&&(1 !=2'b1));assign Kd5dwq2[5]=((((Ts0dwq2 >=32'h35000000)&&(Ts0dwq2 <=32'h3500ffff))
||(((Ts0dwq2 >=32'h36000000)&&(Ts0dwq2 <=32'h3600ffff))&&(0==1'b1)))&&(1 !=2'b1));assign Kd5dwq2[6]=((((Ts0dwq2 >=32'h37000000)&&(Ts0dwq2 <=32'h3700ffff))
||(((Ts0dwq2 >=32'h38000000)&&(Ts0dwq2 <=32'h3800ffff))&&(0==1'b1)))&&(1 !=2'b1));assign Kd5dwq2[7]=((((Ts0dwq2 >=32'h39000000)&&(Ts0dwq2 <=32'h3900ffff))
||(((Ts0dwq2 >=32'h3a000000)&&(Ts0dwq2 <=32'h3a00ffff))&&(0==1'b1)))&&(1 !=2'b1));assign Kd5dwq2[8]=((((Ts0dwq2 >=32'h3b000000)&&(Ts0dwq2 <=32'h3b00ffff))
||(((Ts0dwq2 >=32'h3c000000)&&(Ts0dwq2 <=32'h3c00ffff))&&(0==1'b1)))&&(1 !=2'b1));assign Kd5dwq2[9]=((((Ts0dwq2 >=32'h3d000000)&&(Ts0dwq2 <=32'h3d00ffff))
||(((Ts0dwq2 >=32'h3e000000)&&(Ts0dwq2 <=32'h3e00ffff))&&(0==1'b1)))&&(1 !=2'b1));assign Kd5dwq2[10]=((((Ts0dwq2 >=32'h3f000000)&&(Ts0dwq2 <=32'h3f00ffff))
||(((Ts0dwq2 >=32'h40000000)&&(Ts0dwq2 <=32'h4000ffff))&&(0==1'b1)))&&(1 !=2'b1));assign Kd5dwq2[11]=((((Ts0dwq2 >=32'h41000000)&&(Ts0dwq2 <=32'h4100ffff))
||(((Ts0dwq2 >=32'h42000000)&&(Ts0dwq2 <=32'h4200ffff))&&(0==1'b1)))&&(1 !=2'b1));assign Kd5dwq2[12]=((((Ts0dwq2 >=32'h43000000)&&(Ts0dwq2 <=32'h4300ffff))
||(((Ts0dwq2 >=32'h44000000)&&(Ts0dwq2 <=32'h4400ffff))&&(0==1'b1)))&&(1 !=2'b1));assign Kd5dwq2[13]=((((Ts0dwq2 >=32'h45000000)&&(Ts0dwq2 <=32'h4500ffff))
||(((Ts0dwq2 >=32'h46000000)&&(Ts0dwq2 <=32'h4600ffff))&&(0==1'b1)))&&(1 !=2'b1));assign Kd5dwq2[14]=((((Ts0dwq2 >=32'h47000000)&&(Ts0dwq2 <=32'h4700ffff))
||(((Ts0dwq2 >=32'h48000000)&&(Ts0dwq2 <=32'h4800ffff))&&(0==1'b1)))&&(1 !=2'b1));assign Kd5dwq2[15]=((((Ts0dwq2 >=32'h49000000)&&(Ts0dwq2 <=32'h4900ffff))
||(((Ts0dwq2 >=32'h4a000000)&&(Ts0dwq2 <=32'h4a00ffff))&&(0==1'b1)))&&(1 !=2'b1));assign Xd5dwq2=(Sc5dwq2 ? Ad5dwq2[2:0]: Kd5dwq2[2:0]);
assign Os0dwq2[2:0]=Xd5dwq2;assign Os0dwq2[(2+1)]=Ve0dwq2;always @(Xd5dwq2)begin : Ge5dwq2 Ve0dwq2=1'b1;for(Op0dwq2=0;(Op0dwq2 <=2);Op0dwq2=(Op0dwq2+1))begin 
if(Xd5dwq2[Op0dwq2]==1'b1)begin Ve0dwq2=1'b0;end end end endmodule module A91dwq2(Ve5dwq2,Ud0dwq2,Zd0dwq2,Zs0dwq2,He0dwq2,Kk0dwq2,Rm0dwq2,
Oe0dwq2,Au0dwq2,Pz0dwq2,Wu0dwq2,N01dwq2,M11dwq2,Ym0dwq2,X21dwq2,Mm0dwq2,F51dwq2,Ku0dwq2,Cv0dwq2,Nx0dwq2,Fx0dwq2,F31dwq2);
parameter Df5dwq2=2'b0;parameter Ff5dwq2=2'b1;parameter Hf5dwq2=2'b10;parameter Kf5dwq2=2'b11;output[3:0]Ve5dwq2;input Ud0dwq2;
input Zd0dwq2;input[(3-1):0]Zs0dwq2;input He0dwq2;input[(2-1):0]Kk0dwq2;input[(16-1):0]Rm0dwq2;input[(2-1):0]Oe0dwq2;
input[1:0]Au0dwq2;input[1:0]Ku0dwq2;output[1:0]F51dwq2;input[(4-1):0]Pz0dwq2;input Wu0dwq2;input[1:0]N01dwq2;input M11dwq2;
input[1:0]Ym0dwq2;input X21dwq2;output Mm0dwq2;output[1:0]Cv0dwq2;output Nx0dwq2;output[(4-1):0]Fx0dwq2;output F31dwq2;
reg[3:0]Ve5dwq2;reg[1:0]F51dwq2;reg[1:0]Cv0dwq2;reg[(4-1):0]Fx0dwq2;reg F31dwq2;reg Mf5dwq2;reg Xf5dwq2;reg Hg5dwq2;
reg[1:0]Og5dwq2;reg[1:0]Wg5dwq2;reg[(4-1):0]Gp2dwq2;reg[(4-1):0]Ih5dwq2;reg Uh5dwq2;reg[3:0]Ai5dwq2;reg[3:0]Hi5dwq2;
reg[3:0]Ki5dwq2;reg Oi5dwq2;reg[1:0]Vi5dwq2;reg[1:0]Lj5dwq2;reg[3:0]Yj5dwq2;reg[3:0]Ik5dwq2;reg[3:0]Tk5dwq2;reg[3:0]El5dwq2;
reg[3:0]Pl5dwq2;reg Dm5dwq2;reg[15:0]Jm5dwq2;wire[1:0]Vm5dwq2;wire Gn5dwq2;wire Mn5dwq2;wire Un5dwq2;wire Zn5dwq2;wire Do5dwq2;
wire Lo5dwq2;wire So5dwq2;wire Xo5dwq2;wire Bp5dwq2;wire Op5dwq2;wire Sp5dwq2;wire Gq5dwq2;integer Op0dwq2;integer Qp0dwq2;
integer Yp0dwq2;integer Oq5dwq2;integer Wp0dwq2;integer Qq5dwq2;integer Sq5dwq2;assign Bp5dwq2=(X21dwq2==1'b1);assign Xo5dwq2=((He0dwq2==1'b1)&&((Oe0dwq2==2'b11)||(Oe0dwq2==2'b10)
));assign Sp5dwq2=((Vi5dwq2 !=Cv0dwq2)&&(He0dwq2==1'b1));assign Gq5dwq2=(((Zs0dwq2 > 3'b1)&&(Oe0dwq2==2'b11))&&(Kk0dwq2==2'b0))
;assign Zn5dwq2=(Rm0dwq2[Gp2dwq2]&&(Og5dwq2 !=Df5dwq2));assign Un5dwq2=(Wg5dwq2 !=Df5dwq2);assign Gn5dwq2=((Ai5dwq2==4'b0)&&(Gq5dwq2==1'b0));
assign Mn5dwq2=((Ai5dwq2==4'b1)&&(He0dwq2==1'b1));assign Lo5dwq2=((((((Un5dwq2==1'b1)&&(Kk0dwq2==2'b11))&&(Og5dwq2 !=
Df5dwq2))&&(Dm5dwq2==1'b0))||((Un5dwq2==1'b0)&&((Oe0dwq2 !=2'b1)||(Gn5dwq2==1'b1))))||(Zn5dwq2==1'b1));assign Op5dwq2=(((Kk0dwq2==2'b10)||(Kk0dwq2==2'b11))&&(Wg5dwq2==
Df5dwq2));assign Do5dwq2=(((((Mn5dwq2==1'b1)||(Gn5dwq2==1'b1))&&(Lo5dwq2==1'b1))&&(Sp5dwq2==1'b0))||(Op5dwq2==1'b1));
assign Vm5dwq2={{1 {1'b0}},1'b1};assign So5dwq2=(((He0dwq2==1'b1)&&(Oi5dwq2==1'b1))||(Og5dwq2==Hf5dwq2));assign Nx0dwq2=(Og5dwq2==Ff5dwq2);
assign Mm0dwq2=Hg5dwq2;always @(Au0dwq2 or Ih5dwq2 or Xf5dwq2)begin : Uq5dwq2 Mf5dwq2=1'b0;for(Op0dwq2=0;(Op0dwq2 <=1);Op0dwq2=(Op0dwq2+1))begin 
Mf5dwq2=((((Au0dwq2[Op0dwq2]==1'b1)&&(Ih5dwq2==Op0dwq2))&&(Xf5dwq2==1'b1))|| Mf5dwq2);end end always @(He0dwq2 or Og5dwq2)begin : Kr5dwq2 
if(Og5dwq2==Kf5dwq2)begin Xf5dwq2=1'b0;end else begin Xf5dwq2=He0dwq2;end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Zr5dwq2 
if(Zd0dwq2==1'b0)begin Hg5dwq2 <=1'b0;end else begin if(Xf5dwq2==1'b1)begin Hg5dwq2 <=Mf5dwq2;end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Ls5dwq2 
if(Zd0dwq2==1'b0)begin Uh5dwq2 <=1'b0;end else begin if(Og5dwq2==Kf5dwq2)begin Uh5dwq2 <=1'b1;end else begin Uh5dwq2 <=1'b0;
end end end always @(Kk0dwq2 or Oe0dwq2 or Zs0dwq2 or Hi5dwq2 or Bp5dwq2)begin : Ws5dwq2 if((((((Bp5dwq2==1'b1)||(Kk0dwq2==2'b11))||(Kk0dwq2==2'b10))||(
Oe0dwq2==2'b0))||(Zs0dwq2==3'b0))||(Zs0dwq2==3'b1))begin Ai5dwq2=4'b0;end else begin if(((Zs0dwq2==3'b111)||(Zs0dwq2==3'b110))&&(Oe0dwq2==2'b10))begin 
Ai5dwq2=4'hf;end else begin if(((Zs0dwq2==3'b101)||(Zs0dwq2==3'h4))&&(Oe0dwq2==2'b10))begin Ai5dwq2=4'h7;end else 
begin if(((Zs0dwq2==3'b011)||(Zs0dwq2==3'b010))&&(Oe0dwq2==2'b10))begin Ai5dwq2=4'h3;end else begin if(Hi5dwq2==4'b0)begin 
Ai5dwq2=4'b0;end else begin Ai5dwq2=(Hi5dwq2-4'b1);end end end end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : It5dwq2 
if(Zd0dwq2==1'b0)begin Hi5dwq2 <=4'b0;end else begin if(Xo5dwq2==1'b1)begin Hi5dwq2 <=Ai5dwq2;end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Qt5dwq2 
if(Zd0dwq2==1'b0)begin Vi5dwq2 <={2 {1'b1}};end else begin Vi5dwq2 <=Cv0dwq2;end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Eu5dwq2 
if(Zd0dwq2==1'b0)begin Ki5dwq2 <=4'b0;end else begin if(Xo5dwq2==1'b1)begin Ki5dwq2 <=Ve5dwq2;end end end always @(Zs0dwq2 or Oe0dwq2 or Ki5dwq2)begin : Nu5dwq2 
if(Zs0dwq2 > 3'b1)begin case(Oe0dwq2)2'b10: case(Zs0dwq2[2:1])1: Ve5dwq2=4'h3;2: Ve5dwq2=4'h7;default: Ve5dwq2=4'hf;
endcase 2'b11: Ve5dwq2=(Ki5dwq2-4'b1);2'b0: Ve5dwq2=4'b0;default: Ve5dwq2=Ki5dwq2;endcase end else begin Ve5dwq2=4'b0;
end end always @(Ve5dwq2 or Ku0dwq2 or Fx0dwq2)begin : Av5dwq2 F51dwq2=Ku0dwq2;if(Ve5dwq2 > 4'b1)begin F51dwq2[Fx0dwq2]=1'b1;
end end always @(Ym0dwq2)begin : Ov5dwq2 Jm5dwq2 <=16'b0;Jm5dwq2[1:0]<=Ym0dwq2;end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Fw5dwq2 
if(Zd0dwq2==1'b0)begin Cv0dwq2 <={{1 {1'b0}},1'b1};end else if(Do5dwq2==1'b1)begin if((((Un5dwq2==1'b1)&&(Kk0dwq2==2'b11))||(Bp5dwq2==1'b1))||(Wu0dwq2 
==1'b1))begin Cv0dwq2 <=Vm5dwq2;end else begin if((Zn5dwq2==1'b1)||((Og5dwq2==Hf5dwq2)&&(Kk0dwq2==2'b10)))begin for(Qp0dwq2=0;(Qp0dwq2 <=1);Qp0dwq2=(Qp0dwq2+1))begin 
Cv0dwq2[Qp0dwq2]<=(Gp2dwq2==Qp0dwq2[3:0]);end end else begin if(M11dwq2==1'b1)begin if((Kk0dwq2==2'b10)&&(He0dwq2==1'b0))begin 
for(Qp0dwq2=0;(Qp0dwq2 <=1);Qp0dwq2=(Qp0dwq2+1))begin Cv0dwq2[Qp0dwq2]<=(Gp2dwq2==Qp0dwq2[3:0]);end end else begin 
if(Jm5dwq2[Pz0dwq2]==1'b1)begin Cv0dwq2 <=Vm5dwq2;end else begin for(Qp0dwq2=0;(Qp0dwq2 <=1);Qp0dwq2=(Qp0dwq2+1))begin 
Cv0dwq2[Qp0dwq2]<=(Pz0dwq2==Qp0dwq2[3:0]);end end end end else begin Cv0dwq2 <=N01dwq2;end end end end else begin if(Bp5dwq2==1'b1)begin 
Cv0dwq2 <=Vm5dwq2;end end end always @(Cv0dwq2 or Pz0dwq2)begin : Vw5dwq2 Ih5dwq2=Pz0dwq2;for(Oq5dwq2=0;(Oq5dwq2 <=1);Oq5dwq2=(Oq5dwq2+1))begin 
if(Cv0dwq2[Oq5dwq2]==1'b1)begin Ih5dwq2=Oq5dwq2[3:0];end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Mx5dwq2 
if(Zd0dwq2==1'b0)begin Fx0dwq2 <={4 {1'b0}};end else begin if(He0dwq2==1'b1)begin Fx0dwq2 <=Ih5dwq2;end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Zx5dwq2 
if(Zd0dwq2==1'b0)begin Oi5dwq2 <=1'b0;end else begin if(He0dwq2==1'b1)begin if(Og5dwq2==Df5dwq2)begin Oi5dwq2 <=1'b1;
end else begin Oi5dwq2 <=1'b0;end end end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Ly5dwq2 if(Zd0dwq2==1'b0)begin 
Gp2dwq2 <={4 {1'b0}};end else begin if(So5dwq2==1'b1)begin Gp2dwq2 <=Fx0dwq2;end end end always @(Oe0dwq2 or He0dwq2 or Hg5dwq2)begin : Az5dwq2 
if((((Oe0dwq2==2'b10)||(Oe0dwq2==2'b0))||(Hg5dwq2==1'b1))&&(He0dwq2==1'b1))begin F31dwq2=1'b1;end else begin F31dwq2=1'b0;
end end always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin : Nz5dwq2 if(Zd0dwq2==1'b0)begin Og5dwq2 <=Df5dwq2;end else begin 
Og5dwq2 <=Wg5dwq2;end end always @(Og5dwq2 or He0dwq2 or Mf5dwq2 or Hg5dwq2 or Oe0dwq2 or Uh5dwq2 or  Kk0dwq2 or Ih5dwq2 or Gp2dwq2 or Dm5dwq2)begin : A06dwq2 
case(Og5dwq2)Ff5dwq2: if((He0dwq2==1'b1)&&(Oe0dwq2 !=2'b1))begin if((Mf5dwq2==1'b1)||((Hg5dwq2==1'b1)&&(Uh5dwq2==1'b1)))begin 
Wg5dwq2=Ff5dwq2;end else begin Wg5dwq2=Hf5dwq2;end end else begin if((Kk0dwq2==2'b11)&&(Dm5dwq2==1'b0))begin Wg5dwq2=Kf5dwq2;
end else begin Wg5dwq2=Ff5dwq2;end end Hf5dwq2: if((He0dwq2==1'b1)&&(Oe0dwq2 !=2'b1))begin if((Mf5dwq2==1'b1)||(Kk0dwq2==2'b10))begin 
Wg5dwq2=Ff5dwq2;end else begin Wg5dwq2=Df5dwq2;end end else begin if(Kk0dwq2==2'b11)begin Wg5dwq2=Kf5dwq2;end else begin 
Wg5dwq2=Hf5dwq2;end end Kf5dwq2: if((He0dwq2==1'b1)&&(Ih5dwq2==Gp2dwq2))begin Wg5dwq2=Ff5dwq2;end else begin Wg5dwq2=Kf5dwq2;
end default: if((He0dwq2==1'b1)&&(Mf5dwq2==1'b1))begin Wg5dwq2=Ff5dwq2;end else begin Wg5dwq2=Df5dwq2;end endcase end 
always @(posedge Ud0dwq2 or negedge Zd0dwq2)begin if(Zd0dwq2==1'b0)begin Dm5dwq2 <=1'b0;end else begin if((Og5dwq2==Df5dwq2)&&(Wg5dwq2==Ff5dwq2))begin 
Dm5dwq2 <=1'b1;end else begin if(He0dwq2==1'b1)begin Dm5dwq2 <=1'b0;end end end end endmodule module ahb_wrapper(bus_hbusreq,bus_hgrant,bus_hlock,hsel,hclk,hresetn,pause,
haddr_m1,hburst_m1,hbusreq_m1,hlock_m1,hprot_m1,hsize_m1,htrans_m1,hwdata_m1,hwrite_m1,hgrant_m1,hsel_s1,hready_resp_s1,hresp_s1,hrdata_s1,
hsel_s2,hready_resp_s2,hresp_s2,hrdata_s2,haddr,hburst,hprot,hsize,htrans,hwdata,hwrite,hready,hresp,hrdata,ahbarbint,hmaster,hmaster_data,
hmastlock);output[(4-1):0]hsel;output[1:0]bus_hbusreq;output[1:0]bus_hlock;output[1:0]bus_hgrant;input hclk;input hresetn;
input pause;input[(32-1):0]haddr_m1;input hbusreq_m1;input[(3-1):0]hburst_m1;input hlock_m1;input[(4-1):0]hprot_m1;
input[(3-1):0]hsize_m1;input[(2-1):0]htrans_m1;input[(`L3lkc-1):0]hwdata_m1;input hwrite_m1;output hgrant_m1;input hready_resp_s1;
input[(2-1):0]hresp_s1;input[(`L3lkc-1):0]hrdata_s1;output hsel_s1;input hready_resp_s2;input[(2-1):0]hresp_s2;input[(`L3lkc-1):0]hrdata_s2;
output hsel_s2;output[(32-1):0]haddr;output[(3-1):0]hburst;output[(4-1):0]hprot;output[(3-1):0]hsize;output[(2-1):0]htrans;
output[(`L3lkc-1):0]hwdata;output hwrite;output[(4-1):0]hmaster;output[(4-1):0]hmaster_data;output hmastlock;output ahbarbint;
output hready;output[(2-1):0]hresp;output[(`L3lkc-1):0]hrdata;wire Sc5dwq2;wire[(((1+1)*32)-1):0]Nk1dwq2;wire[(4-1):0]Cm1dwq2;
wire[(32-1):0]Qk0dwq2;wire[(6-1):0]Un1dwq2;wire[(3-1):0]Jn1dwq2;wire[((3*`L3lkc)-1):0]Eo1dwq2;wire[(6-1):0]Xk1dwq2;
wire[(6-1):0]Sl1dwq2;wire[(8-1):0]Il1dwq2;wire[(2-1):0]Ym1dwq2;wire[((2*`L3lkc)-1):0]Nm1dwq2;wire R76dwq2;wire Xv0dwq2;
wire[(`L3lkc-1):0]Vw0dwq2;wire[(2-1):0]Mw0dwq2;wire Ve0dwq2;wire[(2-1):0]Wf0dwq2;wire Ff0dwq2;wire[(`L3lkc-1):0]Hg0dwq2;
wire Z76dwq2;wire J86dwq2;wire[1:1]Xx0dwq2;wire Jy0dwq2;assign Nk1dwq2[(32-1):0]={32 {1'b0}};assign Cm1dwq2[(2-1):0]=2'b0;
assign Nm1dwq2[(`L3lkc-1):0]={`L3lkc {1'b0}};assign Sl1dwq2[(3-1):0]=3'b0;assign Xk1dwq2[(3-1):0]=3'b0;assign Il1dwq2[(4-1):0]=4'hc;
assign Ym1dwq2[0]=1'b0;assign Nk1dwq2[63:32]=haddr_m1;assign Cm1dwq2[3:2]=htrans_m1;assign Xk1dwq2[5:3]=hburst_m1;assign Sl1dwq2[5:3]=hsize_m1;
assign Il1dwq2[7:4]=hprot_m1;assign Ym1dwq2[1]=hwrite_m1;assign Nm1dwq2[((`L3lkc*2)-1):(`L3lkc*1)]=hwdata_m1;assign bus_hbusreq[1]=hbusreq_m1;
assign hgrant_m1=bus_hgrant[1];assign bus_hlock[1]=hlock_m1;assign bus_hbusreq[0]=1'b0;assign bus_hlock[0]=1'b0;assign Jn1dwq2[0]=Xv0dwq2;
assign Un1dwq2[1:0]=Mw0dwq2;assign Eo1dwq2[(`L3lkc-1):0]=Vw0dwq2;assign Jn1dwq2[1]=hready_resp_s1;assign Un1dwq2[3:2]=hresp_s1;
assign Eo1dwq2[((`L3lkc*2)-1):(`L3lkc*1)]=hrdata_s1;assign Jn1dwq2[2]=hready_resp_s2;assign Un1dwq2[5:4]=hresp_s2;assign Eo1dwq2[((`L3lkc*3)-1):(`L3lkc*2)]=hrdata_s2;
assign Ve0dwq2=hsel[(2+1)];assign R76dwq2=hsel[0];assign hsel_s1=hsel[1];assign hsel_s2=hsel[2];assign Qk0dwq2[15:0]={16 {1'b0}};
assign Qk0dwq2[31:16]={16 {1'b0}};assign J86dwq2=((0==1'b1)? Sc5dwq2 : 1'b1);assign Z76dwq2=((1==1'b1)? pause : 1'b0);
Ck1dwq2 V86dwq2(.Ud0dwq2(hclk),.Zd0dwq2(hresetn),.Nk1dwq2(Nk1dwq2),.Xk1dwq2(Xk1dwq2),.Fx0dwq2(hmaster),.Il1dwq2(Il1dwq2),.Sl1dwq2 
(Sl1dwq2),.Cm1dwq2(Cm1dwq2),.Nm1dwq2(Nm1dwq2),.Ym1dwq2(Ym1dwq2),.Hg0dwq2(Hg0dwq2),.Ff0dwq2(Ff0dwq2),.Wf0dwq2(Wf0dwq2),.Jn1dwq2 
(Jn1dwq2),.Un1dwq2(Un1dwq2),.Eo1dwq2(Eo1dwq2),.Os0dwq2(hsel[2:0]),.Bl0dwq2(hmaster_data),.Ts0dwq2(haddr),.Zs0dwq2(hburst),.Po1dwq2 
(hprot),.Gt0dwq2(hsize),.Oe0dwq2(htrans),.Mt0dwq2(hwdata),.Tt0dwq2(hwrite),.Vo1dwq2(hrdata),.He0dwq2(hready),.Kk0dwq2(hresp));
Gc5dwq2 B96dwq2(.Ts0dwq2(haddr),.Sc5dwq2(J86dwq2),.Os0dwq2(hsel));Ds0dwq2 I96dwq2(.Ud0dwq2(hclk),.Zd0dwq2(hresetn),.He0dwq2(hready),
.Kk0dwq2(hresp),.Os0dwq2(R76dwq2),.Ts0dwq2(haddr),.Zs0dwq2(hburst),.Gt0dwq2(hsize),.Oe0dwq2(htrans),.Mt0dwq2(hwdata),.Tt0dwq2(hwrite),
.Au0dwq2(bus_hlock),.Ku0dwq2(bus_hbusreq),.Qk0dwq2(Qk0dwq2),.Bl0dwq2(hmaster_data),.Wu0dwq2(Z76dwq2),.Cv0dwq2(bus_hgrant),.Nv0dwq2 
(ahbarbint),.Xv0dwq2(Xv0dwq2),.Mw0dwq2(Mw0dwq2),.Vw0dwq2(Vw0dwq2),.Fx0dwq2(hmaster),.Nx0dwq2(hmastlock),.Xx0dwq2(Xx0dwq2),.Jy0dwq2 
(Jy0dwq2));Fd0dwq2 O96dwq2(.Ud0dwq2(hclk),.Zd0dwq2(hresetn),.He0dwq2(hready),.Oe0dwq2(htrans),.Ve0dwq2(Ve0dwq2),.Ff0dwq2(Ff0dwq2),.Wf0dwq2 
(Wf0dwq2),.Hg0dwq2(Hg0dwq2));endmodule module V91dwq2(Sa1dwq2,Wa1dwq2,Cb1dwq2,Kb1dwq2,Tb1dwq2,Ym0dwq2,F11dwq2,Yb1dwq2,N31dwq2,H01dwq2,Gc1dwq2);
parameter Up0dwq2=4;parameter Y96dwq2=2;parameter Ga6dwq2=1;parameter Qa6dwq2=0;parameter Bb6dwq2=1;input Sa1dwq2;input Wa1dwq2;
input[(Up0dwq2-1):0]Cb1dwq2;input[(Up0dwq2-1):0]Tb1dwq2;input[(Up0dwq2-1):0]Ym0dwq2;input[((Y96dwq2*Up0dwq2)-1):0]Kb1dwq2;
output F11dwq2;output Yb1dwq2;output N31dwq2;output[(Up0dwq2-1):0]H01dwq2;output[(((Up0dwq2 > 4096)?((Up0dwq2 > 262144)?((Up0dwq2 > 2097152)?((
Up0dwq2 > 8388608)? 24 :((Up0dwq2 > 4194304)? 23 : 22)):((Up0dwq2 > 1048576)? 21 :((Up0dwq2 > 524288)? 20 : 19))):((Up0dwq2 > 32768)?((Up0dwq2 >  
131072)? 18 :((Up0dwq2 > 65536)? 17 : 16)):((Up0dwq2 > 16384)? 15 :((Up0dwq2 > 8192)? 14 : 13)))):((Up0dwq2 > 64)?((Up0dwq2 > 512)?((Up0dwq2 > 
2048)? 12 :((Up0dwq2 > 1024)? 11 : 10)):((Up0dwq2 > 256)? 9 :((Up0dwq2 >  128)? 8 : 7))):((Up0dwq2 > 8)?((Up0dwq2 > 32)? 6 :((Up0dwq2 > 16)? 5 : 4 
)):((Up0dwq2 > 4)? 3 :((Up0dwq2 > 2)? 2 : 1)))))-1):0]Gc1dwq2;integer Wc6dwq2;integer Md6dwq2;reg De6dwq2;reg Pe6dwq2;
reg Bf6dwq2;reg Of6dwq2;reg Ag6dwq2;reg Lg6dwq2;reg[(Up0dwq2-1):0]Wg6dwq2;reg Nh6dwq2;reg Wh6dwq2;reg Gi6dwq2;reg Pi6dwq2;
reg Zi6dwq2;reg Gj6dwq2;reg Ik5dwq2;reg[((Y96dwq2*Up0dwq2)-1):0]Nj6dwq2;integer Fl6dwq2;integer Tl6dwq2;integer Op0dwq2;
integer Nb6dwq2[(Up0dwq2-1):0];integer Ec6dwq2[(Up0dwq2-1):0];integer Ak6dwq2[(Up0dwq2-1):0];integer Qk6dwq2[(Up0dwq2-1):0];
assign H01dwq2=((Wc6dwq2==(-2))? {Up0dwq2 {1'bx}} :(((Md6dwq2==(-1))&&(Bb6dwq2==0))? {Up0dwq2 {1'b0}} :((Bb6dwq2==0)?(1'b1 << Md6dwq2):(1'b1 
<< Wc6dwq2))));assign Gc1dwq2=((Wc6dwq2==(-2))? {((Up0dwq2 > 4096)?((Up0dwq2 > 262144)?((Up0dwq2 > 2097152)?((Up0dwq2 > 8388608)? 24 :((Up0dwq2 > 4194304)? 23 :  
22)):((Up0dwq2 > 1048576)? 21 :((Up0dwq2 > 524288)? 20 : 19))):((Up0dwq2  > 32768)?((Up0dwq2 > 131072)? 18 :((Up0dwq2 > 65536)? 17 : 16)):((Up0dwq2 
> 16384)? 15 :((Up0dwq2 > 8192)? 14 : 13)))):((Up0dwq2 > 64)?((Up0dwq2 >  512)?((Up0dwq2 > 2048)? 12 :((Up0dwq2 > 1024)? 11 : 10)):((Up0dwq2 > 256)
? 9 :((Up0dwq2 > 128)? 8 : 7))):((Up0dwq2 > 8)?((Up0dwq2 > 32)? 6 :((Up0dwq2 > 16)? 5 : 4)):((Up0dwq2 > 4)? 3 :((Up0dwq2 > 2)? 2 : 1))))){1'bx 
}} :(((Wc6dwq2==(-1))&&(Bb6dwq2==1))? {((Up0dwq2 > 4096)?((Up0dwq2 >  262144)?((Up0dwq2 > 2097152)?((Up0dwq2 > 8388608)? 24 :((Up0dwq2 > 4194304 
)? 23 : 22)):((Up0dwq2 > 1048576)? 21 :((Up0dwq2 > 524288)? 20 : 19))):((Up0dwq2 > 32768)?((Up0dwq2 > 131072)? 18 :((Up0dwq2 > 65536)? 17 : 16)):  
((Up0dwq2 > 16384)? 15 :((Up0dwq2 > 8192)? 14 : 13)))):((Up0dwq2 > 64)?((Up0dwq2 > 512)?((Up0dwq2 > 2048)? 12 :((Up0dwq2 > 1024)? 11 : 10)):((
Up0dwq2 > 256)? 9 :((Up0dwq2 > 128)? 8 : 7))):((Up0dwq2 > 8)?((Up0dwq2 >  32)? 6 :((Up0dwq2 > 16)? 5 : 4)):((Up0dwq2 > 4)? 3 :((Up0dwq2 > 2)? 2 :  
1))))){1'b1}} :(((Md6dwq2==(-1))&&(Bb6dwq2==0))? {((Up0dwq2 > 4096)?((Up0dwq2 > 262144)?((Up0dwq2 > 2097152)?((Up0dwq2 > 8388608)? 24 :((
Up0dwq2 > 4194304)? 23 : 22)):((Up0dwq2 > 1048576)? 21 :((Up0dwq2 > 524288)? 20 : 19))):((Up0dwq2 > 32768)?((Up0dwq2 > 131072)? 18 :((Up0dwq2 > 65536 
)? 17 : 16)):((Up0dwq2 > 16384)? 15 :((Up0dwq2 > 8192)? 14 : 13)))):((Up0dwq2 > 64)?((Up0dwq2 > 512)?((Up0dwq2 > 2048)? 12 :((Up0dwq2 > 1024)?  
11 : 10)):((Up0dwq2 > 256)? 9 :((Up0dwq2 > 128)? 8 : 7))):((Up0dwq2 > 8)?((Up0dwq2 > 32)? 6 :((Up0dwq2 > 16)? 5 : 4)):((Up0dwq2 > 4)? 3 :((
Up0dwq2 > 2)? 2 : 1))))){1'b1}} :((Bb6dwq2==0)? Md6dwq2 : Wc6dwq2))));assign Yb1dwq2=((Bb6dwq2==0)? Bf6dwq2 : Pe6dwq2);
assign F11dwq2=((Bb6dwq2==0)? De6dwq2 : Ag6dwq2);assign N31dwq2=((Bb6dwq2==0)? Of6dwq2 : Lg6dwq2);always @(Wc6dwq2 or Pe6dwq2 or Cb1dwq2 or Tb1dwq2 or Ym0dwq2 or Kb1dwq2 or  
Nb6dwq2[0])begin : Nm6dwq2 Pi6dwq2=(^Cb1dwq2);Zi6dwq2=(^Tb1dwq2);Gj6dwq2=(^Ym0dwq2);Ik5dwq2=(^Kb1dwq2);Fl6dwq2=(-1);
Nh6dwq2=1'b0;Wh6dwq2=1'b0;Gi6dwq2=1'b0;for(Op0dwq2=0;(Op0dwq2 < Up0dwq2);Op0dwq2=(Op0dwq2+1))Qk6dwq2[Op0dwq2]=Nb6dwq2[Op0dwq2];
Tl6dwq2=0;Nj6dwq2=Kb1dwq2;for(Op0dwq2=0;(Op0dwq2 < Up0dwq2);Op0dwq2=(Op0dwq2+1))begin Ak6dwq2[Op0dwq2]=Nj6dwq2[(Y96dwq2-1):0];
Nj6dwq2=(Nj6dwq2 >> Y96dwq2);end Wg6dwq2=(Cb1dwq2 &(~Ym0dwq2));if((Wc6dwq2 <(-1))&&(Tb1dwq2 !=={Up0dwq2 {1'b0}}))begin 
Fl6dwq2=(-2);Gi6dwq2=1'bx;Wh6dwq2=1'bx;end else if((Wc6dwq2 >=0)&&(Tb1dwq2[Wc6dwq2]!==1'b0))begin if(Tb1dwq2[Wc6dwq2]===1'b1)begin 
Fl6dwq2=Wc6dwq2;Gi6dwq2=1'b1;Wh6dwq2=1'b1;if(Pe6dwq2===1'b0)begin Tl6dwq2=1;end end else begin Fl6dwq2=(-2);Gi6dwq2=1'bx;
Wh6dwq2=1'bx;Nh6dwq2=1'b0;end end else if(Wg6dwq2 !=={Up0dwq2 {1'b0}})begin if((Pi6dwq2===1'bx)||(Ik5dwq2===1'bx))begin 
Fl6dwq2=(-2);Wh6dwq2=1'bx;Nh6dwq2=1'bx;end else begin for(Op0dwq2=0;(Op0dwq2 < Up0dwq2);Op0dwq2=(Op0dwq2+1))begin 
if(Wg6dwq2[Op0dwq2]===1'b1)begin if((Fl6dwq2 < 0)||((Ak6dwq2[Op0dwq2]< Ak6dwq2[Fl6dwq2])||((Ak6dwq2[Op0dwq2]==Ak6dwq2[Fl6dwq2])&&(Nb6dwq2[Op0dwq2]< Nb6dwq2[Fl6dwq2])))
)begin Fl6dwq2=Op0dwq2;Wh6dwq2=1'b1;end end end Tl6dwq2=1;end end else if(Ga6dwq2==1)begin Fl6dwq2=Qa6dwq2;Nh6dwq2=1'b1;
end else begin Fl6dwq2=(-1);end for(Op0dwq2=0;(Op0dwq2 < Up0dwq2);Op0dwq2=(Op0dwq2+1))begin if(Op0dwq2==Fl6dwq2)begin 
Qk6dwq2[Op0dwq2]=(1 <<(((Up0dwq2 > 4096)?((Up0dwq2 > 262144)?((Up0dwq2 >  2097152)?((Up0dwq2 > 8388608)? 24 :((Up0dwq2 > 4194304)? 23 : 22)):((
Up0dwq2 > 1048576)? 21 :((Up0dwq2 > 524288)? 20 : 19))):((Up0dwq2 > 32768)?((Up0dwq2 > 131072)? 18 :((Up0dwq2 > 65536)? 17 : 16)):((Up0dwq2 > 16384)
? 15 :((Up0dwq2 > 8192)? 14 : 13)))):((Up0dwq2 > 64)?((Up0dwq2 > 512)?((Up0dwq2 > 2048)? 12 :((Up0dwq2 > 1024)? 11 : 10)):((Up0dwq2 > 256)? 9 :((
Up0dwq2 > 128)? 8 : 7))):((Up0dwq2 > 8)?((Up0dwq2 > 32)? 6 :((Up0dwq2 >  16)? 5 : 4)):((Up0dwq2 > 4)? 3 :((Up0dwq2 > 2)? 2 : 1)))))-1));
end else if(Wg6dwq2[Op0dwq2]==1'b1)begin if(Tl6dwq2==1)begin if(Qk6dwq2[Op0dwq2]==0)begin Qk6dwq2[Op0dwq2]=(1 <<(((Up0dwq2 > 4096)?((Up0dwq2 > 262144)?((Up0dwq2 >  
2097152)?((Up0dwq2 > 8388608)? 24 :((Up0dwq2 > 4194304)? 23 : 22)):((Up0dwq2 > 1048576)? 21 :((Up0dwq2 > 524288)? 20 : 19))):((Up0dwq2 > 32768)
?((Up0dwq2 > 131072)? 18 :((Up0dwq2 > 65536)? 17 : 16)):((Up0dwq2 > 16384)? 15 :((Up0dwq2 > 8192)? 14 : 13)))):((Up0dwq2 > 64)?((Up0dwq2 > 512)?((
Up0dwq2 > 2048)? 12 :((Up0dwq2 > 1024)? 11 : 10)):((Up0dwq2 > 256)? 9 :((Up0dwq2 > 128)? 8 : 7))):((Up0dwq2 > 8)?((Up0dwq2 > 32)? 6 :((Up0dwq2 >  
16)? 5 : 4)):((Up0dwq2 > 4)? 3 :((Up0dwq2 > 2)? 2 : 1)))))-1));end else begin Qk6dwq2[Op0dwq2]=(Nb6dwq2[Op0dwq2]-1);end 
end end else begin Qk6dwq2[Op0dwq2]=(1 <<(((Up0dwq2 > 4096)?((Up0dwq2 > 262144)?((Up0dwq2 >  2097152)?((Up0dwq2 > 8388608)? 24 :((Up0dwq2 > 4194304)? 23 : 22)):((
Up0dwq2 > 1048576)? 21 :((Up0dwq2 > 524288)? 20 : 19))):((Up0dwq2 > 32768)?((Up0dwq2 > 131072)? 18 :((Up0dwq2 > 65536)? 17 : 16)):((Up0dwq2 > 16384)
? 15 :((Up0dwq2 > 8192)? 14 : 13)))):((Up0dwq2 > 64)?((Up0dwq2 > 512)?((Up0dwq2 > 2048)? 12 :((Up0dwq2 > 1024)? 11 : 10)):((Up0dwq2 > 256)? 9 :((
Up0dwq2 > 128)? 8 : 7))):((Up0dwq2 > 8)?((Up0dwq2 > 32)? 6 :((Up0dwq2 >  16)? 5 : 4)):((Up0dwq2 > 4)? 3 :((Up0dwq2 > 2)? 2 : 1)))))-1));
end end Md6dwq2=Fl6dwq2;De6dwq2=Nh6dwq2;Bf6dwq2=Wh6dwq2;Of6dwq2=Gi6dwq2;for(Op0dwq2=0;(Op0dwq2 < Up0dwq2);Op0dwq2=(Op0dwq2+1))
Ec6dwq2[Op0dwq2]=Qk6dwq2[Op0dwq2];end always @(posedge Sa1dwq2 or negedge Wa1dwq2)begin : Xm6dwq2 if(Wa1dwq2===1'b0)begin Wc6dwq2 <=(-1);
Ag6dwq2 <=1'b0;Pe6dwq2 <=1'b0;Lg6dwq2 <=1'b0;for(Op0dwq2=0;(Op0dwq2 < Up0dwq2);Op0dwq2=(Op0dwq2+1))Nb6dwq2[Op0dwq2]<=(1 <<(((Up0dwq2 > 4096)?((Up0dwq2 > 262144)?((Up0dwq2 > 
2097152)?((Up0dwq2 > 8388608)? 24 :((Up0dwq2 > 4194304)? 23 : 22)):((Up0dwq2 > 1048576)? 21 :((Up0dwq2 > 524288)? 20 : 19))):((Up0dwq2 > 32768)
?((Up0dwq2 > 131072)? 18 :((Up0dwq2 > 65536)? 17 : 16)):((Up0dwq2 > 16384)? 15 :((Up0dwq2 > 8192)? 14 : 13)))):((Up0dwq2 > 64)?((Up0dwq2 > 512)?((
Up0dwq2 > 2048)? 12 :((Up0dwq2 > 1024)? 11 : 10)):((Up0dwq2 > 256)? 9 :((Up0dwq2 > 128)? 8 : 7))):((Up0dwq2 > 8)?((Up0dwq2 > 32)? 6 :((Up0dwq2 >  
16)? 5 : 4)):((Up0dwq2 > 4)? 3 :((Up0dwq2 > 2)? 2 : 1)))))-1));end else if(Wa1dwq2===1'b1)begin Wc6dwq2 <=Md6dwq2;Ag6dwq2 <=De6dwq2;
Pe6dwq2 <=Bf6dwq2;Lg6dwq2 <=Of6dwq2;for(Op0dwq2=0;(Op0dwq2 < Up0dwq2);Op0dwq2=(Op0dwq2+1))Nb6dwq2[Op0dwq2]<=Ec6dwq2[Op0dwq2];
end else begin Wc6dwq2 <=(-2);Ag6dwq2 <=1'bx;Pe6dwq2 <=1'bx;Lg6dwq2 <=1'bx;for(Op0dwq2=0;(Op0dwq2 < Up0dwq2);Op0dwq2=(Op0dwq2+1))
Nb6dwq2[Op0dwq2]<=(-1);end end initial begin : Gn6dwq2 integer Wn6dwq2;Wn6dwq2=0;if((Up0dwq2 < 2)||(Up0dwq2 > 32))begin 
Wn6dwq2=1;$display("ERROR: %m :\n  Invalid value(%d)for parameter n(legal range: 2 to 32)",Up0dwq2);end if((Y96dwq2 < 1)||(Y96dwq2 > 5))begin 
Wn6dwq2=1;$display("ERROR: %m :\n  Invalid value(%d)for parameter p_width(legal range: 1 to 5)",Y96dwq2);end if((Ga6dwq2 < 0)||(Ga6dwq2 > 1))begin 
Wn6dwq2=1;$display("ERROR: %m :\n  Invalid value(%d)for parameter park_mode(legal range: 0 to 1)",Ga6dwq2);end if((Qa6dwq2 < 0)||(Qa6dwq2 >(Up0dwq2-1)))begin 
Wn6dwq2=1;$display("ERROR: %m :\n  Invalid value(%d)for parameter park_index(legal range: 0 to n-1)",Qa6dwq2);end if((Bb6dwq2 < 0)||(Bb6dwq2 > 1))begin 
Wn6dwq2=1;$display("ERROR: %m :\n  Invalid value(%d)for parameter output_mode(legal range: 0 to 1)",Bb6dwq2);end if(Wn6dwq2==1)begin 
$display("%m :\n  Simulation aborted due to invalid parameter value(s)");$finish;end end always @(Sa1dwq2)begin : Bp6dwq2 if(((Sa1dwq2 !==1'b0)&&(Sa1dwq2 !==1'b1))&&($time > 0))begin 
$display("WARNING: %m :\n  at time=%t,detected unknown value,%b,on clk input.",$time,Sa1dwq2);end end endmodule module Mp1dwq2(Dq1dwq2,Fq1dwq2,Jq1dwq2);
parameter Tp6dwq2=8;parameter Bq6dwq2=2;parameter Lq6dwq2=2;input[(Tp6dwq2-1):0]Dq1dwq2;input[(Bq6dwq2-1):0]Fq1dwq2;
output[(Lq6dwq2-1):0]Jq1dwq2;assign Jq1dwq2=Vq6dwq2(Dq1dwq2,Fq1dwq2);function[(Lq6dwq2-1):0]Vq6dwq2;input[(Tp6dwq2-1):0]Br6dwq2;
input[(Bq6dwq2-1):0]Dr6dwq2;reg[(Tp6dwq2-1):0]Br6dwq2;reg[(Bq6dwq2-1):0]Dr6dwq2;integer Op0dwq2;integer Qp0dwq2;reg[(Lq6dwq2-1):0]Hr6dwq2;
begin for(Op0dwq2=0;(Op0dwq2 < Lq6dwq2);Op0dwq2=(Op0dwq2+1))begin Qp0dwq2=((Dr6dwq2*Lq6dwq2)+Op0dwq2);if(Qp0dwq2 >(Tp6dwq2-1))begin 
Hr6dwq2[Op0dwq2] = 1'b0; end else begin Hr6dwq2[Op0dwq2] = Br6dwq2[Qp0dwq2]; end end Vq6dwq2 = Hr6dwq2; end endfunction endmodule 